
module model_tb #(

  localparam
    CONV2_XB=10, CONV2_KB=5,
    CONV2_XH=8, CONV2_XW=8, CONV2_XC=1, CONV2_YC=32,
    CONV2_KH=5, CONV2_KW=5, CONV2_SH=2, CONV2_SW=2,
    CONV2_YH=CONV2_XH/CONV2_SH, CONV2_YW=CONV2_XW/CONV2_SW,
    CONV2_YB=CONV2_XB+CONV2_KB + $clog2(CONV2_KH*CONV2_KW*CONV2_XC+1),
    CONV2_XD=CONV2_XH*CONV2_XW*CONV2_XC,
    CONV2_KD=CONV2_KH*CONV2_KW*CONV2_XC*CONV2_YC, CONV2_BD=CONV2_YC,
    CONV2_YD=CONV2_YH*CONV2_YW*CONV2_YC,
  localparam
    ACT3_XB=CONV2_YB, ACT3_XBF=9, ACT3_YBQ=11, ACT3_YBI=3, ACT3_D=512, 
    ACT3_NEGATIVE_SLOPE=0,
    ACT3_YB=ACT3_YBQ+(ACT3_NEGATIVE_SLOPE==0),
  localparam
    DENSE5_XD=512, DENSE5_YD=16, DENSE5_KB=7, DENSE5_XB=ACT3_YB,
    DENSE5_YB=DENSE5_XB + DENSE5_KB + $clog2(DENSE5_XD+1),
    DENSE5_KD=DENSE5_XD*DENSE5_YD, DENSE5_BD=DENSE5_YD,
  localparam
    ACT6_XB=DENSE5_YB, ACT6_XBF=13, ACT6_YBQ=13, ACT6_YBI=3, ACT6_D=16, 
    ACT6_NEGATIVE_SLOPE=0,
    ACT6_YB=ACT6_YBQ+(ACT6_NEGATIVE_SLOPE==0),
  localparam
    XD=CONV2_XD, XB=CONV2_XB, 
    YD=ACT6_D, YB=ACT6_YB,
    WEIGHTS_B = 61616);

  wire [WEIGHTS_B-1:0] weights = {  7'd0, 7'd0, 7'd0, 7'd0, 7'd0, 7'd0, 7'd0, 7'd0, 7'd0, 7'd0, 7'd0, 7'd0, 7'd0, 7'd0, 7'd0, 7'd0, 7'd0, -7'd1, -7'd1, -7'd2, 7'd3, -7'd1, 7'd0, 7'd1, -7'd3, 7'd1, 7'd1, 7'd2, 7'd2, 7'd0, 7'd1, -7'd3, 7'd1, 7'd5, -7'd2, 7'd3, 7'd1, 7'd1, 7'd0, 7'd1, 7'd1, -7'd3, 7'd2, 7'd0, -7'd1, 7'd0, 7'd2, -7'd2, -7'd2, 7'd0, -7'd4, -7'd2, 7'd3, 7'd1, -7'd2, 7'd1, 7'd2, 7'd3, 7'd3, 7'd1, 7'd1, 7'd2, -7'd4, 7'd0, 7'd2, 7'd0, -7'd2, 7'd0, 7'd3, -7'd1, -7'd1, 7'd1, 7'd0, 7'd0, -7'd3, -7'd2, 7'd4, -7'd1, 7'd2, 7'd0, 7'd0, -7'd3, 7'd2, 7'd2, -7'd2, 7'd2, -7'd2, 7'd4, 7'd1, -7'd3, -7'd1, 7'd2, 7'd2, 7'd0, 7'd0, 7'd1, 7'd4, 7'd2, 7'd3, -7'd2, 7'd3, 7'd4, -7'd3, -7'd2, -7'd1, -7'd2, -7'd1, 7'd1, 7'd0, 7'd1, 7'd2, 7'd1, 7'd0, -7'd1, 7'd1, -7'd2, -7'd1, -7'd1, 7'd1, -7'd2, 7'd1, 7'd3, -7'd2, 7'd2, 7'd3, -7'd2, 7'd0, 7'd4, 7'd3, -7'd1, -7'd3, -7'd1, -7'd4, -7'd1, 7'd1, -7'd1, -7'd2, 7'd2, 7'd0, -7'd1, -7'd1, 7'd2, 7'd4, 7'd4, 7'd0, 7'd0, 7'd1, -7'd2, 7'd0, 7'd0, 7'd0, -7'd2, 7'd1, 7'd2, -7'd2, 7'd4, -7'd1, 7'd1, -7'd4, -7'd1, 7'd0, -7'd1, 7'd0, -7'd2, 7'd1, 7'd3, 7'd4, -7'd1, 7'd1, 7'd0, -7'd2, 7'd4, -7'd3, 7'd1, -7'd1, 7'd2, -7'd2, 7'd2, -7'd3, 7'd3, 7'd0, 7'd2, 7'd0, -7'd1, 7'd3, 7'd2, 7'd0, -7'd2, -7'd1, -7'd3, -7'd2, 7'd0, 7'd0, 7'd1, 7'd1, 7'd0, 7'd0, -7'd3, -7'd1, 7'd1, 7'd3, 7'd1, -7'd2, -7'd2, 7'd0, -7'd2, -7'd1, 7'd0, 7'd3, 7'd2, 7'd1, -7'd2, -7'd3, 7'd2, 7'd0, 7'd0, 7'd0, -7'd3, 7'd2, 7'd2, -7'd3, -7'd1, -7'd2, 7'd0, 7'd1, 7'd3, -7'd1, 7'd0, 7'd3, 7'd2, -7'd1, 7'd0, 7'd0, 7'd2, 7'd4, 7'd2, 7'd1, 7'd0, 7'd1, -7'd2, 7'd2, -7'd1, 7'd4, -7'd3, 7'd1, 7'd3, 7'd0, -7'd2, 7'd0, -7'd1, 7'd4, -7'd2, -7'd2, 7'd1, 7'd2, -7'd2, 7'd2, 7'd1, 7'd3, 7'd2, -7'd2, 7'd2, -7'd2, 7'd2, -7'd2, 7'd2, -7'd3, 7'd0, 7'd1, 7'd0, -7'd2, 7'd3, -7'd1, -7'd1, -7'd2, -7'd3, -7'd2, 7'd1, 7'd1, 7'd0, -7'd1, 7'd0, 7'd0, 7'd1, 7'd4, -7'd1, 7'd1, -7'd2, 7'd0, 7'd0, -7'd1, 7'd1, 7'd1, 7'd3, 7'd3, 7'd1, 7'd3, 7'd3, 7'd3, 7'd0, -7'd4, -7'd1, -7'd1, -7'd1, 7'd0, -7'd4, 7'd2, 7'd1, -7'd2, -7'd1, 7'd1, 7'd2, 7'd0, 7'd3, 7'd3, -7'd3, -7'd1, 7'd1, 7'd0, 7'd3, 7'd0, 7'd2, 7'd1, -7'd3, -7'd2, -7'd1, 7'd2, -7'd2, 7'd3, 7'd4, 7'd4, 7'd1, -7'd1, -7'd2, 7'd0, 7'd0, 7'd1, -7'd1, 7'd1, 7'd1, 7'd3, 7'd1, 7'd0, -7'd2, 7'd0, -7'd1, 7'd1, 7'd1, 7'd0, 7'd3, -7'd1, -7'd1, 7'd4, 7'd3, 7'd3, 7'd1, 7'd4, 7'd2, 7'd0, 7'd1, 7'd1, 7'd3, -7'd3, 7'd1, 7'd2, -7'd1, -7'd1, 7'd3, 7'd0, -7'd2, 7'd1, 7'd0, -7'd3, -7'd1, -7'd2, 7'd0, -7'd2, -7'd4, 7'd3, -7'd1, -7'd3, 7'd3, 7'd1, -7'd1, -7'd1, 7'd0, 7'd3, 7'd0, 7'd0, -7'd5, 7'd1, -7'd2, -7'd1, -7'd3, 7'd4, -7'd1, 7'd0, -7'd4, -7'd2, -7'd3, 7'd0, -7'd2, -7'd4, -7'd4, 7'd2, -7'd1, 7'd2, 7'd2, 7'd1, 7'd2, -7'd1, 7'd3, 7'd1, 7'd1, -7'd1, 7'd1, 7'd1, 7'd2, 7'd2, 7'd1, 7'd1, 7'd3, 7'd0, 7'd2, 7'd0, 7'd0, -7'd1, 7'd3, -7'd3, 7'd1, 7'd1, 7'd0, 7'd3, 7'd3, -7'd2, 7'd3, -7'd2, 7'd0, 7'd0, 7'd1, 7'd3, -7'd2, -7'd1, 7'd1, 7'd2, 7'd3, 7'd1, -7'd1, 7'd1, -7'd2, -7'd3, 7'd0, -7'd3, 7'd0, 7'd1, 7'd3, 7'd0, 7'd4, 7'd1, 7'd0, -7'd1, 7'd4, -7'd1, -7'd2, 7'd2, -7'd2, -7'd3, 7'd2, 7'd0, -7'd3, -7'd1, 7'd3, 7'd1, -7'd1, -7'd2, -7'd4, -7'd4, 7'd4, 7'd2, 7'd0, -7'd2, 7'd2, 7'd1, -7'd2, 7'd4, 7'd3, 7'd0, 7'd0, 7'd2, 7'd0, 7'd4, 7'd3, -7'd3, 7'd3, -7'd3, -7'd1, 7'd2, -7'd1, -7'd1, 7'd3, -7'd3, 7'd0, 7'd2, 7'd2, -7'd1, -7'd2, 7'd0, 7'd2, -7'd2, -7'd1, -7'd2, -7'd2, 7'd2, 7'd3, 7'd1, 7'd1, 7'd1, -7'd3, 7'd0, -7'd2, 7'd3, -7'd1, 7'd3, 7'd1, 7'd1, -7'd1, 7'd2, 7'd1, -7'd2, -7'd3, -7'd2, 7'd3, -7'd3, 7'd1, 7'd0, 7'd2, -7'd1, 7'd4, -7'd2, 7'd2, 7'd1, 7'd4, 7'd3, 7'd0, -7'd1, 7'd3, 7'd1, -7'd2, -7'd2, -7'd2, -7'd1, -7'd1, 7'd3, 7'd2, 7'd3, -7'd2, 7'd0, -7'd2, 7'd2, -7'd4, 7'd4, 7'd2, -7'd3, 7'd3, -7'd2, 7'd1, 7'd2, 7'd2, 7'd0, -7'd1, 7'd2, -7'd1, -7'd2, 7'd1, 7'd2, -7'd1, -7'd1, 7'd2, -7'd3, 7'd2, -7'd2, 7'd3, -7'd1, 7'd3, 7'd3, 7'd0, 7'd4, 7'd0, -7'd3, -7'd3, 7'd0, 7'd4, 7'd0, -7'd1, -7'd2, 7'd2, 7'd3, 7'd4, -7'd4, 7'd0, 7'd4, -7'd2, -7'd2, -7'd1, -7'd1, 7'd1, 7'd1, -7'd3, 7'd1, -7'd3, 7'd4, -7'd3, 7'd2, -7'd4, 7'd0, 7'd0, 7'd0, 7'd1, -7'd1, -7'd2, 7'd2, -7'd1, 7'd0, -7'd1, -7'd2, 7'd0, 7'd2, 7'd3, 7'd1, -7'd1, -7'd2, 7'd1, -7'd2, 7'd3, 7'd2, 7'd3, 7'd1, 7'd1, 7'd1, -7'd4, 7'd1, 7'd2, -7'd4, 7'd1, 7'd2, 7'd3, 7'd3, 7'd1, 7'd0, 7'd2, -7'd2, -7'd1, -7'd2, -7'd1, 7'd2, 7'd2, 7'd3, 7'd2, -7'd2, 7'd2, 7'd0, 7'd0, -7'd4, 7'd0, -7'd2, 7'd2, -7'd1, 7'd0, 7'd2, 7'd3, 7'd0, 7'd1, -7'd1, -7'd3, -7'd1, -7'd1, 7'd4, 7'd4, 7'd0, -7'd3, 7'd4, -7'd2, -7'd1, -7'd1, -7'd4, 7'd0, 7'd2, 7'd2, 7'd0, 7'd1, 7'd2, 7'd0, -7'd1, -7'd2, 7'd2, 7'd1, -7'd2, -7'd2, -7'd1, 7'd0, -7'd2, 7'd3, 7'd4, 7'd2, -7'd1, -7'd1, 7'd0, 7'd1, -7'd1, 7'd0, -7'd1, 7'd1, 7'd2, 7'd0, 7'd1, -7'd3, 7'd1, -7'd2, 7'd0, 7'd2, 7'd0, -7'd1, 7'd1, -7'd1, 7'd0, 7'd3, 7'd1, -7'd2, 7'd2, -7'd2, 7'd0, -7'd3, -7'd2, 7'd2, 7'd0, -7'd1, 7'd2, 7'd1, 7'd2, -7'd2, 7'd2, 7'd0, -7'd1, 7'd4, -7'd1, 7'd3, -7'd1, 7'd0, 7'd2, -7'd3, -7'd2, -7'd3, 7'd0, -7'd2, 7'd3, 7'd1, -7'd1, -7'd3, -7'd4, -7'd1, 7'd2, 7'd4, 7'd1, 7'd1, 7'd0, 7'd0, 7'd3, -7'd3, -7'd1, -7'd2, -7'd2, -7'd1, -7'd1, -7'd2, -7'd2, 7'd3, -7'd1, 7'd2, 7'd1, -7'd3, -7'd2, 7'd0, 7'd0, 7'd0, -7'd1, 7'd1, 7'd1, -7'd3, 7'd2, -7'd1, 7'd4, -7'd4, -7'd3, 7'd1, 7'd3, 7'd0, 7'd1, 7'd3, 7'd0, -7'd1, 7'd1, -7'd2, 7'd1, -7'd1, -7'd3, -7'd1, 7'd3, -7'd2, 7'd4, 7'd1, 7'd2, 7'd3, 7'd4, 7'd0, 7'd0, 7'd2, -7'd1, 7'd1, 7'd0, 7'd2, -7'd2, 7'd0, 7'd3, -7'd2, 7'd1, 7'd2, -7'd2, -7'd1, -7'd2, 7'd0, 7'd2, 7'd3, -7'd1, 7'd0, -7'd1, -7'd1, 7'd0, 7'd0, -7'd1, 7'd0, -7'd2, 7'd2, 7'd2, -7'd1, 7'd1, 7'd0, -7'd2, -7'd1, 7'd2, 7'd1, 7'd1, -7'd2, 7'd2, -7'd3, 7'd2, 7'd2, 7'd1, -7'd3, -7'd4, -7'd1, 7'd0, 7'd2, 7'd0, -7'd2, 7'd2, 7'd2, 7'd1, -7'd4, -7'd4, -7'd2, 7'd0, -7'd2, 7'd4, -7'd1, 7'd1, -7'd1, -7'd1, 7'd0, -7'd2, -7'd2, 7'd4, -7'd2, 7'd3, -7'd1, 7'd0, -7'd1, -7'd3, 7'd1, -7'd1, 7'd2, -7'd2, 7'd0, -7'd3, -7'd2, -7'd1, 7'd0, -7'd1, 7'd1, -7'd4, -7'd3, -7'd2, -7'd2, 7'd0, 7'd4, 7'd1, 7'd2, -7'd2, -7'd1, 7'd1, 7'd2, -7'd1, -7'd1, 7'd1, -7'd1, -7'd1, -7'd2, 7'd0, 7'd4, 7'd1, 7'd0, 7'd2, 7'd1, -7'd2, 7'd0, 7'd4, -7'd1, -7'd2, 7'd2, -7'd1, -7'd1, 7'd3, 7'd4, -7'd1, -7'd1, 7'd0, -7'd1, -7'd3, -7'd1, 7'd0, 7'd1, -7'd2, 7'd2, 7'd0, 7'd4, 7'd1, 7'd0, 7'd1, 7'd2, -7'd3, 7'd2, 7'd4, 7'd1, -7'd2, -7'd2, -7'd1, 7'd4, -7'd3, -7'd3, 7'd3, -7'd1, -7'd1, 7'd3, 7'd0, 7'd0, -7'd1, -7'd1, 7'd1, -7'd1, 7'd1, -7'd2, -7'd3, 7'd4, 7'd4, 7'd2, 7'd3, 7'd0, 7'd0, -7'd1, -7'd2, -7'd2, -7'd1, -7'd2, -7'd3, 7'd1, -7'd3, 7'd1, 7'd2, 7'd1, 7'd4, 7'd1, 7'd0, 7'd0, -7'd3, -7'd4, 7'd1, 7'd2, -7'd2, -7'd2, 7'd0, 7'd0, 7'd3, -7'd3, 7'd0, -7'd1, 7'd2, 7'd0, 7'd2, -7'd1, 7'd1, 7'd2, -7'd3, -7'd1, 7'd1, 7'd1, 7'd0, -7'd1, 7'd0, 7'd0, 7'd1, 7'd1, 7'd2, -7'd2, -7'd1, 7'd0, -7'd1, -7'd1, 7'd0, 7'd0, -7'd1, -7'd2, 7'd1, 7'd4, -7'd1, 7'd1, -7'd2, -7'd3, -7'd1, 7'd1, -7'd4, -7'd1, 7'd1, 7'd1, 7'd0, -7'd2, 7'd0, 7'd4, 7'd1, 7'd1, 7'd2, -7'd1, 7'd1, -7'd1, 7'd1, -7'd1, -7'd3, -7'd2, -7'd2, 7'd1, 7'd0, 7'd1, 7'd0, -7'd2, 7'd1, 7'd4, -7'd3, 7'd1, -7'd1, 7'd0, 7'd0, 7'd4, -7'd3, 7'd0, 7'd0, -7'd4, 7'd5, -7'd4, 7'd3, 7'd3, -7'd4, 7'd4, -7'd3, -7'd2, 7'd2, -7'd2, 7'd1, 7'd3, 7'd4, 7'd0, 7'd2, 7'd3, 7'd0, 7'd2, 7'd4, 7'd2, -7'd1, 7'd0, -7'd2, 7'd2, 7'd2, -7'd1, 7'd0, 7'd1, -7'd4, 7'd0, 7'd2, -7'd2, -7'd2, 7'd1, -7'd4, -7'd1, -7'd4, -7'd2, -7'd1, 7'd0, 7'd3, 7'd1, 7'd0, -7'd3, 7'd1, 7'd1, 7'd1, -7'd3, 7'd2, 7'd4, 7'd1, 7'd0, 7'd0, -7'd1, -7'd1, -7'd1, -7'd1, -7'd3, 7'd1, 7'd1, 7'd3, 7'd1, 7'd1, 7'd1, -7'd4, 7'd4, 7'd3, -7'd3, -7'd3, 7'd1, 7'd2, -7'd1, -7'd2, 7'd2, 7'd2, 7'd2, 7'd0, 7'd0, 7'd5, 7'd1, -7'd1, 7'd1, 7'd0, 7'd1, -7'd2, 7'd1, -7'd1, -7'd2, 7'd0, -7'd2, -7'd3, -7'd1, -7'd1, -7'd3, -7'd4, -7'd3, -7'd1, 7'd1, -7'd2, -7'd1, 7'd0, -7'd3, 7'd0, 7'd2, -7'd2, -7'd2, 7'd1, 7'd2, -7'd1, -7'd2, 7'd0, 7'd4, -7'd2, 7'd1, -7'd2, 7'd2, -7'd2, 7'd1, 7'd2, -7'd4, -7'd2, -7'd1, -7'd3, 7'd4, -7'd2, 7'd3, 7'd0, 7'd1, -7'd1, 7'd0, 7'd0, 7'd0, -7'd2, 7'd0, -7'd2, 7'd1, 7'd1, -7'd2, 7'd0, 7'd0, 7'd0, 7'd2, 7'd0, -7'd2, -7'd1, 7'd0, -7'd1, 7'd2, 7'd3, -7'd1, -7'd1, -7'd1, 7'd0, -7'd2, -7'd1, -7'd1, 7'd0, 7'd0, 7'd0, 7'd4, -7'd4, -7'd3, 7'd0, 7'd1, -7'd2, -7'd2, -7'd1, 7'd2, 7'd0, 7'd0, 7'd3, 7'd0, 7'd1, -7'd4, 7'd1, -7'd4, 7'd3, -7'd1, -7'd1, 7'd2, -7'd3, -7'd1, 7'd3, 7'd4, -7'd3, 7'd0, 7'd3, -7'd2, 7'd1, 7'd1, 7'd0, -7'd1, -7'd4, -7'd2, -7'd2, -7'd1, 7'd2, 7'd0, 7'd1, 7'd0, -7'd1, 7'd1, -7'd2, 7'd3, -7'd3, -7'd3, 7'd3, 7'd1, 7'd1, -7'd1, 7'd1, 7'd1, 7'd0, 7'd1, 7'd1, -7'd2, 7'd4, 7'd4, -7'd3, 7'd1, 7'd2, -7'd2, 7'd0, -7'd1, 7'd2, 7'd2, 7'd1, 7'd1, -7'd1, 7'd0, 7'd0, 7'd0, 7'd1, 7'd0, -7'd2, 7'd1, 7'd0, 7'd1, 7'd1, 7'd2, 7'd2, 7'd0, -7'd2, 7'd1, -7'd3, -7'd1, 7'd0, 7'd0, 7'd2, 7'd2, -7'd1, 7'd0, 7'd2, -7'd2, 7'd0, -7'd2, 7'd4, 7'd0, 7'd1, -7'd3, -7'd1, 7'd3, 7'd4, 7'd0, -7'd2, 7'd1, -7'd1, -7'd1, 7'd2, 7'd1, 7'd0, 7'd1, -7'd2, 7'd0, -7'd2, 7'd0, 7'd2, 7'd0, -7'd1, -7'd1, -7'd1, 7'd0, 7'd0, -7'd1, -7'd1, 7'd1, -7'd2, 7'd4, 7'd0, 7'd0, -7'd3, 7'd2, -7'd2, 7'd0, 7'd3, 7'd2, 7'd0, -7'd1, 7'd3, -7'd3, 7'd1, 7'd0, -7'd3, 7'd0, 7'd2, 7'd0, -7'd2, 7'd2, 7'd3, 7'd2, 7'd2, 7'd0, 7'd2, 7'd1, -7'd2, -7'd4, -7'd2, 7'd4, -7'd1, -7'd1, 7'd0, 7'd4, 7'd1, -7'd1, -7'd1, 7'd1, 7'd2, -7'd1, -7'd2, 7'd2, 7'd1, -7'd2, 7'd2, 7'd0, 7'd2, 7'd4, -7'd3, 7'd1, -7'd2, 7'd1, 7'd3, 7'd2, -7'd4, 7'd2, 7'd1, 7'd2, -7'd2, 7'd4, -7'd3, 7'd0, 7'd0, -7'd2, 7'd3, 7'd2, -7'd2, 7'd3, 7'd1, 7'd2, -7'd1, -7'd1, -7'd3, -7'd2, 7'd2, -7'd1, -7'd1, -7'd4, -7'd2, 7'd2, 7'd1, 7'd0, -7'd1, -7'd2, 7'd0, -7'd2, -7'd2, -7'd2, 7'd4, 7'd1, 7'd0, 7'd0, 7'd3, 7'd4, 7'd0, -7'd1, 7'd2, -7'd4, 7'd1, 7'd2, -7'd3, 7'd2, -7'd1, 7'd0, 7'd0, 7'd4, 7'd0, -7'd2, 7'd2, -7'd3, 7'd0, 7'd4, 7'd2, 7'd4, -7'd2, -7'd1, 7'd1, -7'd3, 7'd2, 7'd0, -7'd4, -7'd3, -7'd1, -7'd2, -7'd2, -7'd4, 7'd1, -7'd4, -7'd2, -7'd1, 7'd1, -7'd4, 7'd1, 7'd2, 7'd4, -7'd2, -7'd2, -7'd1, 7'd0, -7'd2, 7'd2, 7'd1, 7'd3, -7'd1, 7'd3, 7'd1, 7'd1, -7'd4, -7'd1, -7'd4, 7'd2, 7'd0, -7'd3, 7'd0, 7'd2, 7'd0, 7'd1, 7'd2, -7'd3, -7'd2, 7'd4, 7'd4, 7'd1, -7'd2, -7'd1, 7'd4, 7'd1, -7'd3, -7'd1, -7'd2, -7'd1, -7'd3, 7'd0, 7'd2, 7'd0, -7'd4, 7'd2, 7'd0, 7'd4, -7'd1, -7'd1, -7'd2, -7'd1, 7'd2, 7'd0, -7'd3, -7'd1, 7'd1, 7'd1, -7'd2, -7'd3, 7'd1, -7'd1, 7'd1, -7'd1, -7'd1, -7'd2, 7'd1, -7'd1, 7'd1, 7'd1, -7'd2, -7'd1, 7'd0, 7'd2, 7'd1, -7'd1, 7'd1, 7'd0, -7'd3, -7'd2, -7'd1, 7'd0, 7'd3, 7'd3, -7'd1, 7'd3, -7'd2, 7'd0, 7'd0, -7'd2, 7'd1, -7'd1, 7'd1, -7'd4, 7'd1, -7'd1, 7'd3, 7'd1, -7'd4, -7'd2, -7'd2, 7'd0, 7'd2, 7'd1, -7'd1, -7'd3, 7'd1, -7'd3, 7'd0, -7'd2, 7'd0, 7'd1, 7'd1, 7'd0, 7'd2, -7'd1, -7'd2, -7'd4, -7'd1, 7'd2, 7'd0, 7'd1, 7'd0, -7'd1, 7'd2, -7'd2, -7'd3, -7'd1, -7'd1, 7'd2, -7'd4, -7'd1, -7'd4, 7'd1, -7'd2, 7'd1, 7'd0, -7'd1, 7'd1, 7'd0, -7'd1, -7'd2, 7'd0, 7'd0, 7'd4, -7'd1, -7'd3, -7'd1, -7'd3, 7'd4, 7'd2, 7'd4, 7'd1, -7'd3, 7'd2, -7'd1, 7'd1, -7'd1, -7'd1, -7'd1, -7'd3, 7'd0, 7'd4, -7'd1, -7'd2, 7'd4, 7'd1, 7'd1, -7'd3, 7'd1, 7'd2, 7'd3, -7'd1, 7'd0, 7'd0, 7'd1, -7'd1, -7'd1, 7'd3, 7'd1, -7'd2, 7'd1, 7'd0, -7'd4, -7'd3, 7'd2, 7'd0, -7'd1, 7'd1, -7'd3, 7'd1, -7'd2, -7'd1, 7'd2, 7'd1, -7'd3, -7'd4, -7'd2, 7'd0, 7'd0, 7'd0, 7'd1, -7'd1, -7'd3, 7'd2, -7'd1, -7'd2, 7'd0, 7'd1, 7'd0, 7'd0, -7'd2, 7'd0, 7'd1, 7'd5, -7'd2, 7'd0, 7'd3, 7'd2, -7'd4, 7'd0, -7'd1, 7'd0, 7'd2, 7'd1, 7'd3, -7'd1, -7'd4, -7'd2, 7'd3, 7'd4, 7'd1, -7'd1, -7'd4, 7'd4, -7'd1, 7'd0, -7'd2, -7'd1, -7'd2, -7'd2, 7'd2, -7'd2, 7'd1, -7'd2, -7'd1, 7'd2, 7'd0, 7'd2, 7'd1, 7'd1, 7'd0, -7'd3, 7'd3, 7'd1, -7'd1, -7'd3, -7'd1, 7'd2, 7'd1, -7'd2, -7'd4, 7'd2, 7'd1, 7'd0, 7'd4, -7'd2, -7'd4, 7'd1, 7'd0, 7'd2, 7'd3, 7'd3, 7'd1, 7'd0, 7'd1, -7'd2, 7'd3, 7'd2, -7'd1, -7'd2, -7'd2, -7'd2, 7'd1, -7'd2, 7'd2, 7'd2, -7'd1, 7'd0, -7'd3, 7'd0, 7'd1, 7'd1, 7'd0, 7'd1, 7'd0, 7'd0, -7'd1, -7'd3, 7'd0, 7'd0, 7'd1, -7'd1, -7'd1, 7'd2, 7'd0, -7'd3, -7'd2, 7'd1, -7'd1, 7'd0, -7'd1, 7'd1, -7'd1, -7'd3, -7'd1, 7'd1, 7'd0, 7'd1, 7'd2, 7'd2, 7'd1, 7'd2, -7'd1, 7'd1, -7'd2, 7'd1, 7'd2, 7'd0, -7'd1, -7'd3, -7'd1, 7'd0, 7'd3, 7'd0, 7'd0, 7'd1, 7'd0, 7'd3, -7'd1, 7'd0, 7'd1, 7'd3, -7'd4, 7'd1, 7'd4, 7'd1, -7'd1, 7'd1, 7'd2, 7'd0, -7'd4, -7'd3, -7'd1, 7'd1, -7'd1, 7'd2, 7'd3, 7'd1, 7'd1, 7'd1, -7'd2, 7'd1, -7'd2, -7'd2, 7'd0, -7'd3, 7'd0, -7'd1, -7'd2, 7'd1, 7'd0, 7'd0, 7'd2, 7'd2, -7'd2, 7'd0, -7'd1, -7'd2, 7'd1, 7'd1, -7'd2, -7'd1, 7'd1, -7'd4, 7'd3, 7'd2, -7'd3, 7'd0, 7'd0, 7'd2, -7'd2, 7'd1, -7'd4, 7'd1, -7'd2, -7'd2, -7'd2, -7'd1, 7'd1, -7'd1, -7'd2, 7'd1, 7'd0, 7'd2, -7'd2, 7'd3, -7'd2, -7'd4, 7'd0, 7'd1, -7'd3, -7'd2, -7'd2, 7'd0, -7'd2, -7'd1, 7'd0, 7'd1, -7'd2, 7'd2, -7'd1, 7'd1, 7'd0, 7'd2, 7'd4, 7'd0, 7'd1, 7'd2, 7'd0, -7'd3, -7'd1, -7'd2, 7'd4, 7'd3, -7'd3, -7'd2, 7'd0, 7'd1, 7'd1, 7'd0, -7'd1, 7'd2, -7'd2, -7'd4, -7'd1, 7'd1, -7'd3, 7'd3, -7'd2, 7'd1, -7'd1, -7'd3, 7'd1, 7'd3, 7'd0, 7'd2, 7'd0, 7'd0, 7'd1, 7'd0, -7'd2, 7'd4, -7'd1, -7'd4, 7'd1, -7'd1, -7'd2, 7'd0, 7'd1, -7'd2, -7'd1, 7'd1, 7'd1, 7'd0, 7'd2, 7'd1, -7'd2, 7'd0, -7'd1, 7'd1, 7'd2, -7'd1, -7'd3, -7'd2, -7'd2, -7'd3, 7'd0, 7'd2, 7'd0, -7'd1, -7'd4, 7'd2, 7'd3, 7'd1, 7'd0, 7'd1, -7'd1, -7'd3, 7'd0, -7'd4, 7'd3, 7'd3, 7'd0, -7'd2, 7'd0, -7'd2, 7'd2, 7'd1, 7'd1, 7'd0, -7'd3, 7'd0, -7'd3, 7'd0, -7'd4, 7'd0, -7'd1, -7'd2, -7'd2, -7'd2, 7'd1, 7'd0, 7'd1, 7'd2, 7'd2, -7'd1, 7'd4, 7'd0, 7'd4, 7'd4, 7'd1, -7'd2, 7'd2, -7'd1, 7'd2, 7'd0, 7'd0, 7'd0, -7'd3, -7'd3, 7'd2, -7'd1, 7'd4, -7'd1, -7'd1, 7'd1, 7'd0, 7'd1, -7'd1, -7'd1, -7'd1, 7'd0, 7'd1, -7'd3, -7'd4, -7'd1, -7'd1, 7'd2, -7'd1, -7'd2, 7'd3, -7'd3, 7'd1, 7'd0, 7'd1, 7'd3, 7'd1, -7'd2, 7'd0, -7'd1, -7'd3, 7'd2, 7'd1, -7'd3, 7'd1, 7'd0, 7'd0, 7'd0, 7'd0, -7'd1, 7'd0, 7'd0, -7'd3, 7'd1, 7'd0, -7'd2, -7'd3, 7'd0, 7'd3, 7'd3, -7'd1, 7'd2, -7'd2, 7'd0, 7'd0, 7'd2, 7'd0, 7'd1, 7'd2, 7'd4, -7'd1, 7'd2, -7'd2, -7'd3, 7'd2, -7'd1, 7'd4, 7'd2, 7'd2, -7'd1, -7'd2, 7'd0, -7'd2, 7'd2, -7'd1, 7'd1, 7'd1, -7'd2, -7'd3, 7'd1, 7'd1, 7'd2, -7'd2, 7'd2, -7'd1, -7'd1, -7'd2, 7'd3, -7'd1, -7'd3, -7'd1, -7'd2, 7'd1, 7'd1, -7'd2, 7'd3, -7'd3, -7'd4, -7'd4, -7'd2, 7'd0, 7'd2, -7'd2, 7'd0, -7'd2, -7'd3, 7'd2, -7'd1, 7'd0, 7'd0, 7'd2, 7'd2, 7'd0, 7'd2, 7'd2, 7'd2, 7'd1, 7'd0, -7'd2, 7'd3, 7'd0, 7'd2, 7'd3, 7'd2, -7'd1, -7'd2, 7'd4, 7'd2, -7'd1, -7'd1, 7'd4, 7'd3, 7'd3, 7'd3, -7'd2, -7'd1, 7'd0, -7'd1, -7'd4, -7'd3, 7'd2, -7'd2, 7'd0, 7'd3, -7'd3, 7'd1, 7'd0, -7'd3, 7'd0, 7'd0, 7'd2, 7'd1, -7'd2, 7'd0, 7'd0, 7'd0, 7'd1, 7'd1, 7'd0, 7'd4, -7'd1, 7'd0, 7'd1, -7'd4, -7'd4, -7'd2, 7'd1, 7'd1, 7'd1, 7'd1, 7'd0, 7'd1, 7'd2, 7'd3, 7'd2, 7'd1, 7'd0, 7'd2, -7'd1, 7'd2, 7'd1, 7'd2, -7'd1, 7'd2, -7'd1, -7'd2, 7'd1, 7'd1, 7'd2, 7'd2, 7'd4, -7'd2, -7'd1, 7'd0, 7'd0, 7'd1, 7'd4, -7'd3, -7'd1, 7'd3, 7'd2, 7'd3, -7'd2, -7'd2, -7'd1, 7'd1, 7'd1, -7'd2, 7'd2, 7'd0, 7'd2, 7'd3, -7'd1, -7'd3, 7'd1, -7'd2, -7'd2, -7'd2, 7'd1, 7'd0, 7'd3, 7'd2, -7'd1, 7'd2, 7'd0, 7'd0, 7'd3, 7'd2, -7'd3, -7'd2, 7'd1, 7'd1, 7'd3, 7'd0, 7'd1, -7'd2, -7'd2, 7'd4, -7'd1, 7'd0, -7'd2, 7'd0, 7'd2, 7'd2, -7'd1, -7'd1, 7'd2, -7'd1, 7'd0, 7'd1, -7'd1, -7'd1, 7'd0, 7'd1, 7'd0, -7'd3, 7'd1, -7'd1, -7'd2, 7'd0, 7'd2, 7'd1, -7'd2, -7'd1, 7'd1, -7'd3, -7'd1, -7'd2, 7'd0, 7'd3, -7'd2, -7'd2, 7'd0, 7'd0, 7'd0, -7'd1, -7'd1, 7'd3, -7'd1, 7'd2, 7'd3, -7'd2, -7'd3, -7'd3, 7'd0, 7'd2, 7'd1, -7'd1, -7'd2, -7'd1, 7'd0, 7'd3, 7'd4, 7'd4, -7'd3, -7'd1, -7'd2, 7'd0, -7'd2, -7'd2, 7'd2, 7'd0, -7'd2, 7'd2, -7'd2, -7'd4, -7'd3, 7'd1, -7'd1, 7'd0, 7'd2, -7'd3, 7'd1, 7'd1, -7'd4, 7'd1, 7'd2, -7'd3, 7'd1, -7'd1, 7'd0, 7'd3, -7'd4, 7'd0, 7'd0, 7'd1, -7'd2, 7'd2, 7'd2, 7'd0, 7'd3, 7'd0, 7'd2, -7'd1, 7'd0, -7'd3, 7'd1, -7'd1, 7'd4, -7'd2, 7'd1, -7'd4, -7'd1, -7'd2, 7'd3, -7'd2, -7'd1, 7'd3, 7'd1, 7'd2, 7'd3, 7'd1, -7'd2, 7'd0, 7'd1, -7'd1, -7'd1, 7'd1, 7'd2, -7'd1, 7'd1, 7'd1, -7'd3, 7'd0, 7'd0, 7'd0, 7'd0, 7'd3, -7'd1, -7'd3, -7'd3, 7'd1, 7'd0, 7'd3, -7'd1, 7'd3, 7'd1, -7'd1, 7'd1, 7'd0, 7'd1, -7'd3, 7'd3, 7'd1, 7'd2, 7'd3, 7'd0, 7'd4, 7'd4, 7'd1, 7'd3, 7'd0, 7'd1, -7'd2, -7'd2, 7'd3, -7'd1, -7'd2, -7'd3, -7'd1, -7'd1, 7'd0, 7'd3, -7'd2, -7'd1, -7'd1, -7'd2, 7'd3, -7'd3, -7'd1, -7'd2, 7'd2, -7'd1, 7'd0, 7'd2, -7'd1, 7'd0, -7'd2, 7'd0, 7'd0, 7'd1, -7'd1, -7'd4, 7'd4, 7'd0, -7'd3, -7'd1, -7'd3, -7'd3, -7'd4, 7'd1, 7'd2, -7'd1, -7'd2, -7'd3, 7'd4, -7'd1, -7'd2, 7'd4, 7'd0, 7'd0, -7'd3, -7'd2, -7'd3, 7'd3, 7'd2, 7'd2, -7'd3, -7'd5, -7'd1, 7'd0, -7'd2, -7'd1, 7'd1, 7'd1, 7'd0, -7'd1, -7'd1, 7'd0, 7'd1, 7'd0, 7'd2, -7'd1, 7'd3, -7'd1, -7'd1, -7'd3, -7'd3, -7'd1, 7'd0, 7'd2, 7'd2, -7'd1, -7'd1, -7'd1, 7'd0, 7'd2, -7'd2, 7'd0, -7'd1, -7'd1, 7'd2, 7'd1, 7'd1, 7'd0, 7'd2, -7'd2, 7'd2, -7'd1, 7'd0, -7'd2, -7'd3, -7'd1, 7'd1, 7'd1, -7'd2, 7'd3, -7'd1, 7'd0, 7'd1, -7'd4, 7'd2, -7'd1, 7'd3, -7'd2, 7'd0, -7'd1, 7'd2, -7'd2, 7'd3, 7'd3, -7'd2, -7'd2, 7'd2, -7'd1, 7'd0, -7'd1, -7'd3, -7'd2, 7'd0, 7'd3, -7'd2, 7'd1, -7'd3, -7'd1, 7'd2, 7'd0, 7'd2, 7'd2, -7'd2, 7'd0, 7'd3, 7'd3, -7'd1, 7'd0, -7'd1, 7'd1, -7'd2, -7'd2, -7'd3, -7'd2, 7'd1, 7'd0, 7'd2, -7'd2, 7'd1, 7'd0, 7'd2, -7'd2, 7'd0, 7'd2, 7'd4, 7'd0, 7'd2, 7'd0, 7'd3, 7'd0, -7'd3, 7'd0, 7'd3, -7'd1, 7'd0, 7'd4, -7'd1, 7'd3, -7'd1, 7'd2, 7'd0, 7'd3, 7'd1, -7'd1, 7'd1, 7'd1, 7'd3, 7'd3, -7'd3, -7'd2, -7'd1, 7'd1, 7'd0, 7'd2, -7'd1, 7'd0, -7'd3, -7'd1, 7'd4, 7'd0, 7'd0, 7'd5, 7'd1, -7'd3, 7'd3, 7'd1, 7'd0, -7'd1, 7'd1, -7'd3, -7'd2, -7'd4, -7'd4, 7'd3, 7'd3, 7'd1, -7'd3, 7'd0, -7'd2, -7'd2, 7'd2, -7'd2, 7'd4, 7'd0, 7'd2, 7'd0, 7'd4, -7'd2, 7'd1, 7'd3, 7'd0, -7'd1, 7'd0, -7'd1, -7'd1, 7'd1, 7'd0, 7'd3, 7'd1, -7'd1, -7'd2, -7'd1, -7'd1, 7'd4, -7'd1, -7'd2, -7'd2, 7'd0, 7'd0, -7'd2, 7'd1, -7'd1, -7'd3, 7'd2, 7'd0, 7'd2, 7'd2, 7'd3, -7'd1, -7'd1, -7'd2, 7'd2, -7'd3, -7'd1, -7'd1, -7'd1, 7'd0, 7'd2, 7'd3, -7'd1, -7'd3, -7'd1, -7'd3, -7'd2, 7'd0, -7'd3, -7'd2, 7'd0, 7'd0, -7'd2, 7'd1, 7'd3, 7'd0, 7'd2, 7'd0, -7'd3, 7'd1, 7'd1, 7'd1, 7'd1, 7'd0, -7'd3, -7'd2, -7'd1, 7'd4, 7'd0, 7'd0, -7'd3, -7'd1, 7'd2, 7'd1, -7'd1, 7'd2, -7'd3, 7'd2, -7'd1, 7'd2, 7'd2, 7'd0, 7'd0, 7'd0, 7'd1, -7'd2, 7'd3, -7'd1, 7'd2, -7'd3, 7'd1, 7'd1, -7'd1, 7'd2, 7'd2, 7'd4, 7'd1, -7'd1, 7'd1, 7'd3, -7'd2, 7'd2, 7'd1, 7'd1, -7'd1, 7'd1, -7'd2, 7'd1, 7'd1, 7'd2, 7'd1, 7'd3, 7'd0, 7'd1, 7'd2, -7'd3, 7'd3, -7'd1, 7'd1, 7'd2, -7'd1, 7'd1, 7'd2, -7'd1, 7'd0, -7'd3, 7'd0, 7'd1, -7'd2, -7'd1, -7'd4, 7'd3, 7'd4, 7'd0, 7'd1, -7'd1, 7'd2, 7'd1, 7'd0, 7'd1, -7'd2, -7'd2, 7'd2, 7'd2, 7'd2, 7'd1, 7'd3, -7'd2, -7'd2, 7'd0, -7'd3, 7'd1, 7'd0, 7'd1, -7'd1, -7'd4, -7'd3, 7'd3, 7'd1, 7'd2, -7'd2, -7'd1, 7'd2, 7'd1, -7'd3, 7'd0, 7'd2, 7'd0, 7'd2, 7'd1, -7'd1, 7'd0, 7'd0, 7'd0, 7'd0, 7'd2, 7'd2, 7'd0, 7'd2, 7'd0, -7'd1, 7'd1, 7'd1, 7'd4, -7'd2, 7'd1, -7'd3, -7'd1, 7'd1, 7'd0, -7'd2, 7'd1, 7'd0, 7'd1, 7'd1, 7'd2, 7'd1, 7'd3, 7'd2, 7'd1, -7'd2, 7'd3, -7'd2, -7'd3, 7'd3, 7'd1, 7'd1, 7'd2, -7'd4, 7'd1, -7'd1, 7'd1, 7'd3, 7'd2, 7'd2, -7'd3, -7'd1, 7'd0, 7'd0, -7'd1, 7'd2, 7'd1, -7'd4, -7'd3, -7'd3, 7'd1, -7'd1, 7'd1, -7'd1, -7'd3, -7'd2, -7'd1, 7'd0, 7'd1, -7'd4, -7'd1, -7'd1, -7'd3, 7'd0, -7'd1, 7'd0, 7'd2, 7'd1, -7'd1, -7'd1, 7'd1, 7'd3, 7'd0, 7'd0, 7'd0, -7'd1, -7'd3, 7'd3, -7'd2, 7'd1, 7'd2, 7'd2, 7'd3, -7'd1, 7'd2, 7'd0, 7'd0, 7'd0, -7'd2, 7'd1, 7'd0, -7'd2, 7'd4, 7'd3, -7'd2, 7'd1, -7'd1, -7'd2, 7'd0, -7'd3, 7'd1, 7'd0, 7'd1, -7'd1, 7'd2, -7'd2, 7'd3, -7'd2, -7'd1, -7'd2, 7'd0, -7'd1, 7'd3, -7'd4, -7'd1, 7'd3, 7'd3, 7'd2, 7'd1, -7'd1, 7'd1, 7'd0, -7'd2, 7'd4, 7'd1, 7'd1, -7'd1, 7'd2, -7'd1, -7'd5, -7'd1, -7'd2, -7'd3, 7'd2, 7'd1, 7'd0, -7'd2, 7'd1, 7'd2, 7'd4, 7'd4, 7'd2, 7'd0, -7'd3, 7'd0, -7'd3, -7'd1, -7'd4, -7'd3, -7'd1, 7'd1, 7'd2, 7'd0, -7'd4, 7'd0, 7'd1, -7'd1, 7'd0, 7'd0, 7'd1, 7'd1, 7'd2, 7'd4, 7'd4, -7'd2, 7'd2, -7'd2, -7'd4, 7'd2, 7'd2, 7'd0, 7'd2, 7'd1, 7'd0, -7'd2, -7'd3, -7'd1, -7'd1, 7'd3, 7'd3, 7'd1, 7'd2, 7'd0, -7'd2, -7'd4, 7'd0, -7'd3, 7'd0, 7'd1, 7'd1, 7'd1, 7'd2, -7'd4, -7'd2, 7'd0, 7'd2, 7'd1, 7'd1, -7'd1, 7'd0, -7'd1, -7'd4, 7'd0, 7'd3, -7'd1, -7'd2, 7'd4, 7'd1, -7'd2, 7'd1, 7'd0, 7'd3, 7'd0, 7'd0, -7'd1, -7'd4, -7'd1, 7'd3, 7'd0, 7'd0, -7'd3, -7'd2, -7'd2, 7'd0, 7'd0, 7'd1, 7'd0, -7'd1, 7'd1, 7'd3, 7'd1, 7'd0, 7'd2, 7'd0, 7'd4, 7'd0, -7'd1, -7'd2, 7'd2, -7'd1, 7'd2, -7'd3, 7'd1, -7'd1, -7'd1, 7'd2, 7'd2, 7'd2, -7'd1, -7'd2, 7'd0, 7'd1, 7'd0, 7'd1, -7'd2, -7'd3, 7'd1, -7'd1, 7'd0, 7'd1, -7'd1, -7'd1, -7'd3, 7'd1, -7'd1, 7'd4, -7'd1, 7'd4, -7'd2, 7'd1, 7'd0, 7'd0, -7'd4, 7'd2, 7'd1, -7'd1, 7'd2, -7'd1, -7'd2, -7'd4, 7'd2, -7'd1, 7'd4, -7'd4, 7'd0, 7'd0, 7'd4, 7'd0, 7'd1, 7'd1, 7'd1, 7'd1, -7'd2, -7'd4, 7'd0, -7'd2, -7'd3, -7'd3, -7'd2, 7'd3, -7'd4, 7'd1, 7'd1, 7'd2, 7'd4, 7'd0, 7'd3, -7'd1, 7'd1, 7'd1, 7'd3, -7'd4, -7'd1, -7'd2, -7'd2, 7'd0, -7'd2, 7'd2, 7'd0, 7'd4, -7'd2, 7'd0, -7'd4, 7'd0, -7'd2, 7'd0, 7'd3, 7'd0, -7'd2, 7'd1, 7'd0, -7'd2, -7'd3, 7'd0, 7'd0, -7'd2, -7'd1, -7'd2, -7'd1, 7'd4, 7'd0, -7'd1, 7'd2, -7'd2, 7'd0, -7'd1, -7'd3, -7'd2, 7'd1, 7'd4, 7'd3, -7'd2, 7'd1, -7'd4, 7'd2, 7'd1, 7'd0, -7'd1, 7'd2, 7'd1, -7'd3, 7'd2, 7'd3, -7'd1, 7'd2, 7'd3, -7'd2, 7'd0, -7'd1, -7'd1, 7'd1, -7'd4, -7'd2, -7'd1, 7'd0, 7'd2, 7'd0, -7'd2, 7'd0, 7'd1, 7'd1, 7'd3, 7'd0, 7'd1, 7'd3, 7'd0, -7'd1, 7'd2, 7'd1, -7'd1, -7'd2, -7'd2, 7'd0, 7'd1, 7'd1, -7'd3, -7'd2, 7'd0, -7'd3, -7'd3, 7'd3, 7'd1, -7'd3, 7'd0, 7'd1, 7'd4, -7'd2, 7'd0, 7'd2, 7'd0, 7'd1, 7'd2, 7'd1, -7'd1, 7'd4, 7'd3, 7'd2, 7'd4, 7'd1, -7'd1, 7'd3, 7'd1, -7'd2, 7'd3, 7'd1, 7'd0, -7'd1, -7'd2, 7'd2, 7'd1, 7'd2, 7'd0, 7'd0, 7'd3, 7'd2, 7'd2, 7'd3, 7'd0, 7'd0, -7'd3, 7'd2, 7'd1, 7'd1, 7'd2, -7'd3, 7'd1, 7'd0, -7'd1, -7'd2, 7'd1, -7'd1, 7'd4, 7'd2, 7'd2, -7'd3, -7'd4, -7'd1, 7'd2, 7'd2, -7'd2, -7'd1, 7'd0, 7'd1, 7'd0, -7'd1, 7'd0, 7'd0, 7'd2, 7'd1, 7'd1, -7'd3, 7'd1, 7'd0, -7'd2, 7'd1, 7'd0, -7'd4, 7'd4, 7'd0, 7'd1, -7'd3, -7'd1, -7'd1, -7'd2, -7'd3, 7'd2, 7'd4, 7'd1, 7'd2, -7'd1, 7'd1, 7'd0, 7'd2, -7'd2, -7'd2, -7'd2, 7'd3, 7'd1, 7'd2, -7'd2, 7'd2, 7'd0, 7'd0, 7'd4, 7'd1, -7'd1, 7'd1, -7'd1, -7'd3, 7'd0, -7'd2, 7'd2, 7'd1, 7'd2, -7'd3, 7'd3, -7'd2, 7'd1, 7'd3, -7'd2, 7'd2, 7'd3, -7'd3, -7'd1, -7'd1, 7'd0, -7'd1, -7'd1, -7'd1, -7'd2, 7'd0, 7'd1, -7'd1, 7'd2, 7'd0, -7'd1, 7'd1, -7'd1, -7'd2, 7'd0, 7'd4, 7'd1, 7'd2, 7'd1, -7'd1, 7'd0, 7'd2, -7'd4, 7'd2, -7'd1, 7'd0, -7'd3, 7'd1, 7'd1, 7'd1, -7'd3, 7'd1, 7'd1, 7'd2, 7'd0, 7'd2, -7'd1, 7'd0, 7'd2, 7'd2, 7'd4, 7'd0, 7'd3, -7'd1, 7'd0, 7'd0, 7'd2, -7'd2, 7'd4, -7'd1, 7'd1, -7'd1, -7'd1, 7'd0, 7'd1, -7'd1, 7'd2, 7'd2, -7'd2, 7'd3, -7'd1, 7'd2, -7'd1, -7'd2, 7'd1, 7'd2, -7'd1, -7'd1, 7'd2, 7'd4, 7'd4, 7'd3, -7'd3, 7'd2, 7'd1, 7'd1, 7'd2, 7'd0, -7'd2, -7'd4, 7'd2, 7'd0, -7'd1, 7'd1, -7'd2, 7'd3, -7'd1, 7'd1, 7'd0, 7'd2, 7'd2, -7'd3, -7'd4, 7'd1, -7'd1, 7'd1, -7'd3, 7'd0, 7'd0, 7'd0, 7'd4, 7'd3, 7'd0, 7'd0, 7'd0, 7'd1, -7'd1, -7'd2, -7'd1, 7'd4, 7'd0, -7'd2, -7'd1, -7'd1, -7'd3, 7'd1, 7'd0, 7'd0, 7'd0, 7'd1, 7'd3, -7'd1, 7'd1, 7'd0, 7'd0, -7'd2, -7'd2, 7'd1, 7'd0, -7'd1, -7'd3, 7'd0, -7'd1, -7'd1, 7'd1, -7'd1, 7'd0, -7'd4, 7'd1, -7'd4, -7'd2, 7'd3, 7'd1, 7'd2, -7'd2, 7'd2, 7'd3, -7'd2, 7'd1, 7'd4, -7'd3, 7'd3, 7'd1, -7'd4, 7'd2, -7'd3, -7'd1, -7'd1, -7'd2, 7'd3, 7'd4, 7'd3, 7'd1, -7'd1, -7'd1, 7'd3, 7'd2, -7'd1, 7'd0, 7'd2, 7'd1, -7'd4, -7'd3, 7'd1, 7'd2, 7'd1, -7'd1, 7'd0, -7'd3, 7'd4, -7'd1, -7'd4, 7'd2, 7'd0, 7'd1, 7'd4, 7'd0, 7'd0, 7'd3, 7'd3, 7'd0, -7'd1, 7'd0, 7'd3, 7'd0, -7'd2, -7'd3, 7'd2, 7'd1, -7'd2, -7'd2, 7'd3, -7'd2, 7'd2, 7'd1, -7'd1, -7'd2, 7'd4, -7'd1, -7'd2, 7'd0, 7'd0, 7'd3, -7'd1, -7'd2, 7'd3, 7'd0, 7'd1, 7'd2, 7'd3, 7'd2, 7'd4, 7'd0, -7'd2, 7'd0, 7'd0, 7'd0, 7'd1, -7'd2, 7'd1, 7'd0, -7'd3, 7'd2, -7'd1, 7'd3, -7'd3, 7'd0, 7'd1, 7'd4, 7'd0, -7'd2, 7'd1, 7'd3, -7'd2, 7'd2, 7'd1, -7'd3, -7'd2, 7'd3, 7'd2, 7'd2, 7'd0, 7'd0, -7'd3, -7'd3, 7'd2, -7'd3, 7'd2, -7'd1, -7'd2, 7'd0, -7'd1, 7'd2, -7'd1, -7'd3, -7'd1, -7'd1, 7'd0, 7'd0, -7'd3, 7'd2, 7'd2, 7'd1, -7'd2, -7'd3, 7'd4, 7'd2, -7'd1, 7'd0, 7'd1, -7'd1, 7'd3, 7'd0, -7'd1, 7'd2, 7'd1, -7'd2, 7'd0, -7'd1, -7'd5, 7'd2, 7'd0, 7'd2, 7'd1, 7'd0, 7'd0, -7'd2, 7'd1, 7'd0, -7'd3, 7'd1, 7'd1, -7'd2, -7'd2, -7'd4, 7'd3, 7'd1, 7'd0, -7'd1, -7'd1, 7'd2, -7'd2, 7'd3, 7'd3, -7'd2, -7'd1, 7'd4, 7'd3, 7'd0, 7'd1, 7'd1, 7'd0, 7'd0, 7'd0, 7'd2, -7'd2, 7'd2, -7'd1, 7'd4, -7'd2, 7'd1, 7'd1, -7'd1, 7'd0, 7'd0, -7'd3, -7'd1, 7'd0, -7'd2, -7'd1, -7'd1, -7'd1, 7'd0, 7'd2, -7'd1, -7'd1, 7'd2, 7'd1, -7'd2, -7'd1, 7'd2, 7'd2, 7'd3, 7'd3, 7'd2, 7'd0, 7'd0, 7'd1, 7'd0, 7'd1, 7'd3, -7'd1, 7'd2, -7'd4, -7'd3, 7'd0, -7'd1, 7'd1, -7'd1, 7'd0, 7'd0, 7'd2, -7'd1, 7'd3, 7'd0, 7'd1, 7'd1, 7'd2, -7'd2, -7'd4, 7'd0, 7'd0, 7'd0, -7'd1, 7'd3, -7'd3, -7'd1, 7'd2, -7'd2, 7'd1, 7'd0, -7'd1, 7'd1, -7'd4, 7'd4, 7'd1, -7'd2, -7'd1, 7'd2, 7'd1, -7'd2, 7'd1, 7'd1, -7'd1, 7'd0, 7'd4, -7'd1, -7'd2, 7'd1, -7'd3, -7'd2, 7'd1, -7'd1, 7'd1, 7'd0, -7'd1, 7'd0, 7'd1, 7'd1, 7'd0, 7'd0, 7'd1, -7'd1, 7'd2, 7'd3, -7'd1, 7'd0, 7'd0, 7'd1, 7'd0, -7'd1, -7'd2, -7'd3, 7'd0, 7'd1, 7'd1, 7'd1, 7'd0, -7'd1, 7'd3, 7'd0, -7'd3, 7'd0, 7'd0, -7'd3, -7'd2, 7'd3, 7'd4, 7'd0, 7'd0, 7'd4, -7'd4, 7'd2, 7'd1, -7'd3, -7'd4, 7'd1, 7'd1, -7'd2, -7'd2, 7'd3, 7'd1, -7'd2, 7'd0, -7'd1, 7'd2, 7'd1, 7'd4, -7'd3, 7'd0, -7'd1, 7'd0, -7'd4, -7'd3, -7'd2, 7'd3, 7'd2, 7'd1, 7'd3, -7'd1, -7'd1, -7'd4, -7'd1, -7'd2, 7'd0, -7'd2, 7'd0, -7'd3, 7'd2, -7'd2, -7'd1, -7'd2, 7'd1, -7'd1, 7'd0, 7'd4, -7'd4, -7'd2, 7'd2, 7'd4, 7'd2, 7'd4, 7'd0, 7'd2, 7'd3, 7'd2, 7'd0, 7'd2, -7'd2, -7'd2, 7'd3, 7'd1, -7'd1, 7'd3, 7'd0, -7'd1, -7'd2, 7'd1, 7'd1, 7'd1, 7'd0, 7'd3, -7'd1, -7'd1, -7'd3, -7'd1, -7'd4, 7'd1, 7'd0, 7'd3, -7'd3, -7'd2, 7'd0, 7'd0, -7'd2, 7'd4, -7'd3, -7'd3, 7'd0, -7'd4, -7'd3, -7'd2, -7'd2, 7'd2, 7'd2, 7'd4, 7'd2, 7'd0, 7'd0, -7'd1, 7'd2, 7'd2, 7'd1, 7'd2, 7'd0, 7'd2, -7'd1, -7'd2, 7'd1, 7'd2, -7'd1, 7'd1, 7'd1, 7'd3, 7'd3, -7'd1, 7'd2, 7'd0, 7'd1, -7'd1, 7'd0, -7'd1, 7'd1, -7'd4, 7'd0, 7'd3, -7'd4, -7'd3, 7'd4, 7'd1, -7'd1, 7'd0, -7'd1, 7'd2, 7'd1, 7'd0, 7'd0, -7'd1, -7'd1, -7'd2, -7'd1, -7'd1, -7'd1, 7'd2, -7'd1, 7'd2, -7'd1, -7'd1, -7'd1, 7'd2, -7'd1, -7'd4, -7'd4, 7'd3, -7'd4, 7'd1, -7'd1, 7'd2, -7'd3, 7'd0, 7'd1, 7'd1, 7'd3, 7'd2, 7'd2, 7'd0, 7'd0, 7'd2, 7'd1, 7'd0, -7'd3, -7'd1, 7'd2, 7'd4, 7'd4, 7'd3, -7'd1, -7'd1, 7'd0, 7'd0, -7'd1, -7'd2, 7'd2, 7'd0, 7'd0, 7'd0, -7'd2, 7'd0, -7'd3, 7'd2, 7'd1, -7'd1, 7'd1, 7'd2, -7'd3, 7'd1, -7'd1, 7'd3, -7'd3, 7'd2, -7'd1, -7'd2, 7'd2, 7'd2, -7'd1, 7'd1, -7'd2, 7'd0, -7'd1, -7'd1, -7'd1, 7'd4, -7'd3, 7'd2, 7'd2, 7'd0, 7'd2, 7'd2, 7'd0, 7'd2, -7'd1, 7'd4, -7'd1, -7'd3, 7'd2, -7'd2, 7'd1, 7'd2, 7'd3, -7'd2, 7'd3, 7'd4, 7'd3, -7'd1, -7'd2, -7'd4, 7'd3, 7'd1, 7'd3, -7'd3, 7'd0, -7'd3, -7'd4, -7'd3, -7'd2, -7'd1, 7'd1, 7'd1, 7'd0, 7'd0, -7'd2, -7'd1, 7'd1, 7'd0, -7'd3, 7'd1, -7'd3, -7'd1, -7'd1, -7'd2, 7'd1, 7'd1, -7'd2, 7'd2, 7'd1, 7'd2, 7'd2, -7'd4, 7'd2, 7'd5, 7'd0, 7'd3, 7'd2, 7'd4, 7'd2, 7'd1, 7'd3, -7'd1, 7'd1, 7'd2, -7'd2, 7'd1, -7'd2, -7'd2, -7'd1, 7'd2, 7'd1, 7'd1, 7'd0, -7'd2, 7'd0, 7'd0, 7'd0, 7'd2, 7'd4, 7'd0, 7'd1, 7'd3, 7'd3, -7'd1, 7'd0, -7'd2, -7'd2, -7'd2, 7'd0, 7'd0, 7'd1, -7'd2, -7'd2, -7'd1, -7'd3, 7'd2, -7'd1, -7'd2, -7'd1, 7'd0, 7'd2, 7'd1, -7'd4, 7'd2, 7'd1, -7'd1, 7'd1, -7'd2, -7'd2, 7'd2, -7'd4, -7'd1, -7'd2, -7'd3, -7'd1, 7'd1, 7'd3, -7'd2, -7'd1, -7'd1, -7'd5, 7'd2, 7'd0, -7'd1, -7'd3, 7'd0, -7'd1, -7'd2, -7'd4, 7'd1, -7'd3, 7'd2, 7'd1, -7'd4, -7'd1, -7'd2, 7'd3, -7'd1, -7'd2, 7'd3, -7'd1, -7'd2, -7'd3, -7'd1, 7'd2, 7'd1, 7'd0, 7'd3, 7'd4, 7'd0, 7'd0, 7'd0, 7'd2, -7'd1, 7'd1, 7'd4, -7'd3, 7'd0, 7'd3, -7'd1, -7'd2, 7'd4, -7'd1, 7'd1, 7'd2, 7'd0, 7'd2, -7'd2, -7'd3, -7'd3, 7'd3, -7'd2, 7'd0, 7'd1, -7'd2, -7'd1, -7'd3, -7'd2, 7'd3, 7'd3, -7'd2, 7'd1, 7'd0, -7'd2, -7'd1, -7'd1, 7'd1, 7'd1, -7'd1, 7'd3, 7'd0, 7'd2, -7'd3, 7'd0, -7'd2, 7'd2, 7'd2, -7'd2, -7'd3, -7'd2, -7'd2, 7'd2, 7'd1, 7'd2, 7'd2, -7'd2, -7'd1, 7'd1, 7'd2, 7'd2, -7'd1, 7'd3, 7'd2, 7'd3, -7'd3, 7'd0, -7'd1, -7'd2, 7'd2, 7'd3, -7'd1, 7'd2, 7'd2, 7'd4, -7'd1, 7'd1, 7'd1, 7'd0, -7'd1, 7'd2, 7'd3, -7'd1, 7'd2, 7'd0, 7'd2, 7'd2, -7'd2, -7'd2, 7'd0, -7'd1, -7'd2, 7'd1, 7'd0, -7'd1, 7'd2, 7'd2, -7'd1, -7'd4, 7'd2, 7'd0, 7'd0, -7'd1, -7'd2, 7'd4, -7'd3, 7'd3, -7'd2, 7'd0, 7'd1, -7'd3, 7'd2, -7'd2, 7'd2, -7'd2, 7'd2, -7'd1, -7'd2, 7'd2, -7'd1, 7'd0, -7'd3, 7'd3, 7'd2, 7'd1, -7'd1, 7'd2, 7'd2, 7'd2, -7'd4, 7'd4, 7'd1, -7'd2, -7'd1, 7'd3, 7'd2, -7'd2, -7'd1, 7'd0, 7'd0, 7'd1, -7'd2, 7'd1, 7'd3, -7'd3, 7'd4, -7'd4, 7'd3, 7'd0, 7'd0, -7'd4, -7'd1, 7'd0, -7'd2, -7'd1, 7'd0, -7'd1, 7'd0, 7'd2, 7'd2, 7'd0, 7'd2, -7'd3, -7'd3, -7'd1, 7'd1, -7'd4, 7'd0, 7'd0, -7'd1, -7'd2, 7'd1, 7'd0, -7'd4, 7'd0, 7'd0, -7'd1, 7'd4, 7'd0, 7'd0, 7'd1, 7'd1, 7'd1, 7'd3, 7'd1, 7'd1, 7'd2, 7'd1, 7'd2, 7'd2, -7'd2, -7'd1, 7'd2, -7'd2, 7'd1, 7'd0, -7'd1, 7'd2, -7'd2, -7'd3, -7'd2, 7'd3, 7'd0, -7'd2, 7'd2, 7'd1, 7'd0, -7'd1, 7'd0, -7'd1, 7'd0, -7'd3, 7'd1, -7'd3, 7'd3, 7'd3, -7'd1, 7'd3, 7'd3, 7'd0, -7'd2, 7'd4, 7'd0, 7'd0, -7'd3, 7'd1, -7'd2, -7'd3, -7'd4, 7'd2, -7'd5, 7'd2, 7'd3, -7'd1, -7'd1, -7'd2, 7'd1, 7'd4, 7'd0, 7'd1, -7'd1, -7'd1, 7'd1, 7'd0, 7'd0, -7'd1, -7'd1, -7'd3, 7'd3, -7'd1, 7'd3, 7'd1, -7'd1, -7'd2, 7'd1, 7'd0, 7'd1, 7'd0, -7'd1, 7'd3, -7'd3, 7'd0, -7'd2, 7'd0, 7'd1, 7'd3, -7'd1, 7'd0, 7'd1, 7'd0, 7'd0, -7'd1, 7'd2, 7'd1, 7'd1, -7'd1, -7'd2, 7'd2, 7'd2, -7'd1, 7'd1, -7'd3, 7'd1, -7'd1, 7'd0, -7'd3, 7'd0, -7'd1, -7'd3, -7'd1, 7'd1, 7'd3, -7'd3, 7'd4, 7'd0, -7'd1, 7'd2, -7'd2, 7'd2, 7'd2, 7'd2, 7'd3, -7'd2, -7'd1, -7'd1, -7'd3, 7'd1, 7'd0, 7'd0, 7'd2, 7'd3, 7'd2, 7'd4, 7'd3, 7'd3, -7'd2, 7'd4, 7'd1, -7'd1, 7'd2, 7'd3, -7'd2, -7'd2, 7'd1, -7'd1, 7'd0, 7'd2, -7'd2, 7'd2, 7'd0, -7'd3, -7'd2, -7'd1, 7'd0, 7'd1, -7'd3, 7'd0, -7'd2, -7'd1, -7'd1, -7'd3, 7'd1, -7'd2, 7'd2, 7'd0, 7'd0, -7'd1, 7'd2, -7'd2, -7'd3, -7'd3, 7'd1, -7'd4, -7'd1, -7'd2, -7'd3, 7'd0, 7'd0, -7'd3, 7'd0, 7'd3, 7'd1, -7'd2, -7'd1, -7'd4, -7'd2, 7'd1, -7'd2, 7'd3, 7'd2, 7'd4, -7'd3, 7'd0, 7'd3, 7'd0, -7'd1, -7'd2, 7'd2, 7'd0, 7'd4, 7'd3, -7'd1, 7'd0, 7'd1, 7'd0, -7'd1, 7'd0, 7'd1, 7'd0, 7'd2, 7'd0, 7'd0, -7'd2, 7'd0, 7'd1, 7'd1, -7'd1, 7'd2, 7'd1, 7'd1, -7'd1, 7'd0, -7'd3, 7'd3, 7'd0, 7'd2, -7'd3, -7'd3, 7'd3, -7'd2, 7'd2, 7'd3, 7'd3, 7'd0, 7'd2, 7'd2, 7'd0, -7'd3, -7'd3, -7'd3, 7'd0, -7'd2, 7'd1, 7'd4, 7'd0, 7'd0, 7'd1, 7'd1, 7'd2, -7'd3, -7'd1, -7'd1, 7'd2, -7'd2, -7'd1, -7'd1, -7'd2, -7'd1, -7'd3, -7'd1, 7'd1, -7'd2, 7'd1, -7'd3, 7'd3, 7'd3, -7'd2, 7'd2, 7'd4, -7'd1, -7'd2, 7'd1, -7'd2, 7'd2, 7'd1, 7'd1, -7'd5, 7'd3, -7'd2, -7'd3, 7'd0, 7'd1, -7'd1, 7'd4, -7'd3, -7'd2, 7'd1, 7'd0, -7'd1, -7'd1, -7'd4, 7'd3, 7'd3, -7'd1, -7'd4, 7'd2, 7'd0, 7'd1, -7'd3, 7'd0, -7'd2, 7'd3, -7'd1, 7'd0, 7'd4, 7'd1, 7'd1, -7'd3, 7'd1, -7'd2, -7'd2, 7'd0, -7'd2, 7'd0, -7'd1, 7'd1, 7'd1, 7'd1, 7'd3, 7'd3, -7'd3, -7'd3, -7'd1, 7'd2, -7'd2, 7'd0, -7'd2, -7'd3, 7'd4, 7'd3, 7'd0, 7'd2, 7'd2, -7'd2, -7'd2, -7'd1, -7'd2, -7'd1, 7'd2, 7'd1, 7'd1, 7'd1, 7'd1, 7'd2, 7'd0, 7'd1, -7'd2, 7'd1, 7'd1, 7'd1, 7'd2, -7'd1, -7'd2, -7'd2, 7'd2, 7'd4, 7'd0, -7'd1, -7'd3, 7'd0, 7'd0, -7'd2, 7'd2, -7'd4, 7'd1, 7'd1, -7'd2, -7'd1, -7'd2, 7'd4, 7'd2, 7'd2, 7'd0, 7'd2, 7'd2, 7'd0, -7'd1, -7'd2, -7'd1, 7'd1, 7'd1, -7'd2, 7'd4, -7'd2, 7'd1, 7'd2, 7'd2, -7'd1, 7'd0, -7'd4, 7'd3, 7'd2, -7'd2, -7'd1, 7'd1, -7'd1, -7'd4, -7'd4, 7'd1, 7'd3, 7'd4, -7'd1, 7'd4, 7'd2, 7'd0, -7'd3, 7'd1, 7'd2, -7'd1, -7'd2, -7'd2, 7'd0, 7'd1, 7'd0, -7'd2, 7'd0, 7'd0, 7'd0, -7'd3, -7'd2, 7'd2, -7'd2, -7'd2, 7'd0, -7'd2, 7'd0, 7'd1, 7'd0, 7'd1, 7'd3, 7'd0, 7'd3, 7'd2, 7'd0, -7'd1, 7'd0, 7'd1, -7'd2, 7'd1, 7'd2, 7'd4, -7'd1, 7'd2, 7'd0, 7'd3, 7'd3, 7'd2, -7'd1, 7'd0, -7'd1, -7'd1, 7'd0, 7'd2, -7'd2, 7'd0, -7'd2, 7'd1, -7'd3, 7'd1, 7'd4, -7'd3, 7'd2, 7'd3, 7'd0, 7'd2, 7'd2, 7'd2, 7'd2, -7'd2, 7'd1, 7'd1, 7'd4, 7'd2, 7'd3, 7'd2, 7'd0, 7'd4, -7'd1, -7'd1, 7'd1, 7'd1, -7'd4, 7'd4, -7'd1, 7'd1, -7'd2, 7'd3, -7'd2, -7'd1, 7'd0, 7'd3, -7'd2, -7'd1, -7'd1, 7'd3, 7'd0, 7'd2, 7'd0, 7'd1, 7'd0, -7'd1, -7'd3, 7'd3, -7'd1, 7'd0, 7'd1, -7'd4, -7'd2, -7'd2, -7'd1, 7'd1, 7'd1, 7'd1, 7'd1, -7'd2, -7'd1, 7'd0, 7'd0, -7'd1, -7'd1, -7'd2, 7'd3, 7'd0, -7'd1, -7'd2, 7'd2, -7'd2, 7'd0, -7'd5, -7'd1, 7'd1, 7'd3, -7'd2, -7'd4, -7'd1, -7'd3, -7'd1, -7'd1, 7'd3, -7'd2, -7'd2, 7'd1, 7'd1, -7'd3, -7'd4, -7'd2, 7'd2, -7'd1, 7'd1, -7'd2, 7'd0, 7'd0, 7'd0, 7'd3, -7'd2, -7'd1, -7'd4, 7'd1, 7'd2, -7'd1, -7'd3, -7'd1, -7'd1, 7'd0, 7'd2, 7'd1, -7'd2, 7'd3, 7'd1, -7'd1, 7'd5, 7'd2, 7'd1, 7'd1, -7'd1, 7'd2, 7'd2, -7'd2, 7'd1, -7'd2, 7'd0, -7'd2, 7'd2, 7'd4, 7'd1, 7'd0, 7'd0, 7'd0, -7'd1, 7'd1, 7'd0, -7'd4, -7'd2, 7'd3, -7'd3, 7'd3, 7'd1, 7'd1, -7'd1, -7'd2, 7'd0, -7'd3, 7'd2, -7'd1, 7'd1, -7'd1, 7'd3, -7'd1, 7'd1, 7'd1, -7'd3, -7'd4, -7'd3, 7'd1, -7'd3, -7'd1, 7'd0, 7'd2, -7'd4, 7'd1, -7'd1, 7'd4, 7'd0, -7'd1, 7'd0, -7'd1, 7'd3, 7'd1, 7'd1, 7'd4, -7'd3, 7'd0, -7'd1, 7'd3, 7'd0, 7'd0, 7'd1, -7'd1, -7'd2, -7'd1, 7'd0, -7'd3, 7'd2, -7'd3, -7'd1, -7'd1, 7'd2, 7'd0, -7'd4, 7'd2, 7'd1, 7'd0, -7'd1, 7'd4, 7'd2, 7'd3, -7'd1, 7'd3, 7'd2, 7'd3, -7'd2, 7'd2, 7'd3, -7'd1, 7'd1, -7'd1, -7'd1, -7'd1, 7'd1, -7'd2, 7'd2, -7'd3, -7'd3, 7'd3, -7'd1, 7'd4, 7'd5, 7'd2, -7'd2, 7'd0, -7'd2, 7'd0, 7'd4, -7'd1, 7'd1, 7'd2, 7'd3, 7'd2, 7'd0, 7'd2, 7'd0, 7'd0, -7'd1, 7'd1, 7'd1, -7'd1, -7'd1, 7'd2, -7'd1, 7'd3, 7'd3, -7'd2, -7'd4, -7'd3, -7'd2, 7'd3, 7'd2, 7'd4, -7'd1, -7'd1, -7'd2, -7'd3, 7'd3, -7'd1, 7'd0, -7'd2, -7'd1, 7'd0, 7'd0, -7'd4, 7'd2, -7'd1, 7'd1, 7'd3, 7'd2, -7'd3, 7'd0, 7'd4, 7'd1, 7'd1, 7'd2, 7'd0, -7'd2, 7'd0, 7'd1, 7'd0, 7'd3, 7'd2, 7'd0, -7'd2, -7'd2, -7'd1, -7'd2, 7'd3, 7'd0, -7'd3, -7'd1, -7'd1, -7'd1, -7'd1, 7'd3, 7'd0, 7'd0, 7'd2, -7'd1, 7'd0, -7'd2, 7'd2, 7'd0, 7'd1, 7'd0, 7'd0, 7'd1, 7'd2, 7'd1, -7'd1, 7'd0, -7'd2, 7'd2, 7'd3, -7'd2, 7'd0, -7'd1, 7'd2, 7'd0, -7'd3, -7'd2, 7'd1, 7'd0, 7'd0, 7'd0, -7'd1, -7'd1, 7'd2, -7'd4, -7'd2, -7'd4, 7'd5, 7'd2, 7'd1, 7'd0, 7'd1, -7'd4, 7'd3, 7'd1, 7'd0, 7'd3, 7'd2, 7'd2, 7'd0, 7'd1, -7'd2, 7'd1, -7'd4, -7'd2, -7'd3, 7'd1, -7'd1, -7'd1, -7'd1, 7'd2, -7'd1, 7'd1, -7'd1, -7'd1, -7'd1, 7'd3, -7'd1, -7'd3, 7'd2, 7'd2, 7'd2, 7'd1, -7'd2, 7'd2, 7'd1, 7'd0, 7'd0, 7'd4, -7'd3, -7'd1, -7'd3, 7'd2, 7'd3, -7'd1, -7'd1, 7'd0, -7'd1, 7'd0, 7'd3, 7'd4, 7'd4, -7'd4, -7'd2, -7'd3, -7'd3, 7'd1, -7'd1, 7'd0, -7'd1, 7'd1, -7'd2, 7'd1, 7'd2, 7'd0, -7'd1, 7'd1, -7'd2, 7'd1, -7'd2, 7'd2, -7'd3, 7'd2, -7'd2, -7'd1, -7'd2, -7'd2, -7'd1, -7'd2, -7'd4, -7'd2, -7'd4, 7'd1, -7'd1, -7'd3, -7'd3, -7'd2, 7'd1, 7'd3, 7'd4, -7'd1, -7'd2, -7'd2, 7'd0, -7'd2, -7'd2, -7'd2, -7'd1, 7'd1, 7'd1, -7'd3, 7'd3, 7'd1, 7'd1, 7'd2, -7'd2, -7'd3, 7'd0, -7'd1, 7'd4, 7'd0, 7'd0, -7'd2, 7'd1, -7'd3, -7'd1, -7'd3, 7'd0, 7'd3, 7'd0, 7'd0, 7'd1, 7'd4, 7'd1, -7'd2, 7'd0, -7'd1, 7'd0, 7'd0, -7'd4, 7'd0, -7'd2, -7'd3, -7'd1, 7'd0, 7'd2, 7'd2, 7'd3, -7'd2, 7'd1, -7'd1, 7'd3, 7'd0, 7'd1, -7'd1, 7'd0, -7'd2, 7'd0, -7'd1, -7'd2, 7'd1, -7'd1, -7'd2, 7'd0, 7'd1, 7'd0, 7'd4, 7'd1, -7'd1, 7'd0, -7'd2, -7'd2, 7'd2, -7'd2, 7'd0, 7'd2, -7'd3, 7'd0, 7'd0, 7'd2, -7'd2, -7'd1, -7'd2, 7'd0, 7'd3, 7'd1, 7'd1, 7'd1, 7'd2, -7'd1, 7'd4, -7'd1, 7'd3, -7'd4, 7'd2, 7'd0, -7'd2, 7'd1, 7'd4, -7'd1, -7'd3, 7'd1, 7'd0, 7'd1, -7'd2, 7'd0, 7'd0, 7'd3, 7'd0, -7'd3, -7'd3, 7'd1, 7'd4, -7'd2, 7'd0, 7'd1, -7'd3, 7'd0, 7'd1, -7'd2, -7'd2, 7'd0, -7'd2, -7'd1, 7'd1, -7'd2, 7'd0, -7'd2, -7'd4, 7'd1, 7'd1, -7'd2, 7'd0, -7'd1, -7'd2, 7'd2, 7'd0, 7'd0, -7'd3, 7'd0, 7'd0, 7'd3, -7'd1, -7'd1, -7'd2, -7'd3, -7'd2, 7'd2, 7'd1, 7'd2, -7'd2, 7'd1, -7'd1, 7'd2, 7'd0, 7'd2, -7'd2, -7'd4, -7'd2, -7'd3, 7'd3, -7'd3, -7'd1, 7'd1, -7'd1, 7'd2, 7'd3, -7'd1, -7'd2, -7'd2, -7'd2, -7'd3, 7'd4, 7'd2, 7'd0, 7'd0, 7'd0, -7'd3, -7'd4, -7'd1, -7'd1, 7'd0, 7'd3, 7'd0, -7'd1, 7'd1, -7'd2, -7'd3, -7'd2, -7'd3, -7'd2, 7'd1, 7'd1, -7'd4, -7'd2, 7'd2, -7'd4, -7'd1, 7'd1, 7'd0, -7'd3, 7'd2, 7'd0, 7'd1, -7'd5, 7'd1, 7'd3, -7'd1, 7'd4, 7'd1, -7'd2, 7'd2, 7'd4, -7'd1, -7'd1, 7'd1, 7'd0, 7'd4, 7'd0, -7'd2, -7'd3, 7'd0, 7'd1, -7'd4, -7'd1, -7'd4, 7'd3, 7'd0, -7'd3, 7'd1, -7'd2, 7'd2, 7'd1, 7'd1, -7'd3, -7'd3, -7'd3, 7'd3, 7'd0, 7'd2, -7'd1, -7'd2, 7'd1, -7'd2, -7'd2, 7'd1, 7'd0, -7'd3, 7'd0, -7'd3, 7'd3, 7'd1, 7'd0, -7'd4, 7'd1, -7'd1, 7'd0, 7'd0, 7'd0, -7'd2, -7'd1, 7'd3, 7'd0, -7'd3, -7'd2, -7'd1, 7'd1, 7'd1, -7'd2, -7'd2, 7'd3, -7'd2, 7'd4, 7'd1, 7'd1, -7'd1, -7'd1, 7'd3, 7'd0, -7'd1, 7'd4, -7'd1, -7'd1, 7'd2, -7'd3, 7'd1, 7'd2, -7'd2, -7'd1, 7'd1, -7'd2, 7'd1, 7'd1, -7'd2, -7'd3, 7'd0, 7'd0, 7'd1, -7'd1, 7'd2, -7'd1, -7'd3, 7'd2, -7'd1, 7'd2, -7'd1, -7'd2, -7'd1, 7'd0, 7'd3, -7'd3, -7'd1, -7'd1, 7'd2, -7'd1, -7'd4, 7'd0, -7'd1, 7'd2, 7'd1, 7'd1, -7'd2, 7'd1, -7'd2, 7'd3, -7'd1, 7'd1, -7'd2, -7'd3, 7'd3, 7'd3, 7'd0, 7'd3, 7'd1, -7'd2, -7'd3, 7'd1, 7'd0, 7'd0, 7'd0, 7'd0, -7'd2, 7'd0, -7'd1, 7'd0, 7'd4, -7'd2, 7'd1, -7'd1, 7'd0, 7'd3, -7'd1, -7'd1, -7'd1, 7'd2, -7'd2, -7'd1, 7'd0, 7'd1, -7'd3, -7'd3, 7'd2, -7'd1, 7'd1, -7'd1, 7'd0, 7'd1, -7'd1, 7'd1, -7'd1, -7'd2, 7'd0, 7'd0, -7'd1, 7'd0, 7'd3, 7'd0, 7'd1, 7'd4, 7'd2, -7'd3, -7'd1, 7'd0, -7'd2, -7'd4, 7'd0, 7'd0, -7'd2, 7'd2, -7'd1, 7'd2, 7'd0, -7'd1, -7'd2, 7'd3, 7'd3, 7'd1, 7'd2, -7'd3, 7'd0, 7'd1, 7'd0, 7'd1, 7'd1, 7'd3, -7'd2, -7'd1, 7'd1, -7'd1, 7'd1, -7'd3, -7'd3, 7'd0, 7'd2, 7'd4, 7'd2, 7'd2, -7'd1, 7'd0, 7'd4, -7'd2, 7'd0, 7'd2, 7'd1, 7'd2, -7'd4, 7'd1, -7'd2, -7'd2, 7'd1, -7'd1, -7'd1, 7'd0, -7'd4, 7'd2, -7'd2, -7'd2, 7'd0, -7'd3, -7'd1, -7'd1, 7'd1, 7'd0, 7'd3, 7'd0, 7'd1, 7'd2, 7'd1, -7'd2, -7'd3, 7'd0, 7'd1, 7'd3, -7'd1, 7'd3, -7'd2, 7'd1, -7'd4, 7'd0, 7'd0, -7'd2, 7'd2, -7'd2, 7'd0, 7'd0, -7'd2, -7'd3, -7'd1, 7'd0, 7'd0, 7'd0, 7'd3, 7'd0, 7'd1, 7'd1, 7'd3, -7'd2, 7'd1, -7'd2, -7'd3, 7'd2, -7'd3, -7'd2, 7'd3, 7'd2, 7'd0, -7'd1, 7'd3, 7'd3, -7'd4, -7'd1, 7'd1, 7'd2, 7'd1, 7'd2, 7'd2, -7'd1, -7'd1, 7'd4, -7'd2, 7'd3, 7'd2, -7'd1, -7'd1, 7'd1, 7'd0, 7'd0, -7'd1, 7'd2, 7'd0, 7'd0, 7'd1, -7'd1, 7'd0, 7'd1, -7'd3, 7'd1, 7'd3, 7'd2, 7'd0, 7'd1, 7'd4, 7'd2, -7'd1, 7'd1, 7'd4, -7'd1, 7'd2, 7'd3, 7'd1, -7'd1, 7'd3, 7'd2, 7'd2, 7'd3, -7'd2, 7'd2, 7'd0, 7'd2, 7'd3, 7'd1, -7'd1, -7'd2, -7'd4, -7'd4, 7'd0, 7'd3, 7'd2, 7'd1, 7'd0, -7'd2, 7'd3, -7'd2, 7'd1, 7'd0, 7'd0, -7'd1, -7'd1, 7'd1, -7'd1, 7'd0, 7'd1, -7'd2, 7'd2, 7'd0, 7'd1, 7'd0, 7'd2, 7'd1, 7'd0, 7'd3, 7'd1, 7'd0, 7'd0, 7'd2, 7'd0, -7'd1, 7'd3, -7'd1, 7'd0, 7'd1, -7'd4, -7'd1, -7'd1, -7'd2, 7'd0, -7'd2, 7'd0, 7'd0, 7'd1, 7'd2, 7'd0, 7'd4, 7'd0, -7'd1, -7'd2, 7'd1, 7'd2, 7'd2, 7'd3, 7'd1, -7'd1, -7'd2, 7'd0, 7'd1, -7'd3, -7'd2, 7'd1, -7'd1, 7'd1, 7'd1, -7'd1, 7'd0, 7'd1, 7'd1, -7'd2, -7'd1, 7'd1, 7'd1, 7'd0, 7'd3, 7'd0, 7'd1, 7'd4, 7'd2, 7'd2, 7'd0, 7'd0, 7'd4, -7'd4, 7'd1, -7'd2, 7'd2, 7'd0, 7'd3, 7'd0, 7'd1, 7'd3, 7'd3, -7'd2, 7'd2, 7'd1, -7'd2, -7'd1, -7'd3, 7'd1, 7'd0, 7'd1, -7'd4, 7'd4, 7'd1, 7'd0, 7'd0, -7'd2, -7'd3, 7'd0, -7'd1, 7'd1, -7'd1, 7'd3, -7'd4, -7'd3, -7'd1, -7'd3, -7'd2, -7'd3, -7'd2, 7'd1, -7'd1, 7'd3, -7'd1, 7'd1, 7'd1, 7'd0, 7'd2, 7'd1, 7'd3, 7'd4, 7'd0, 7'd4, -7'd1, 7'd3, -7'd2, 7'd1, 7'd0, 7'd0, -7'd1, -7'd1, 7'd3, 7'd0, -7'd2, -7'd2, -7'd2, 7'd1, -7'd2, 7'd0, 7'd0, 7'd0, -7'd3, 7'd0, 7'd0, 7'd0, 7'd3, 7'd3, -7'd3, -7'd1, -7'd4, -7'd1, 7'd1, 7'd0, 7'd1, -7'd2, 7'd1, 7'd1, -7'd2, 7'd0, 7'd0, 7'd0, 7'd5, 7'd1, -7'd1, 7'd3, -7'd1, -7'd4, 7'd2, 7'd0, -7'd2, 7'd0, 7'd0, -7'd1, -7'd1, 7'd4, 7'd1, 7'd1, 7'd4, -7'd2, 7'd2, -7'd2, -7'd3, 7'd1, 7'd2, 7'd2, -7'd4, 7'd4, -7'd2, -7'd2, -7'd1, 7'd2, -7'd4, -7'd2, 7'd1, -7'd2, -7'd2, 7'd3, -7'd2, 7'd0, 7'd1, -7'd1, 7'd2, -7'd3, 7'd2, 7'd0, -7'd3, -7'd1, -7'd1, 7'd1, 7'd2, -7'd2, -7'd1, 7'd0, 7'd2, -7'd1, 7'd0, 7'd1, 7'd2, 7'd2, 7'd2, 7'd2, 7'd1, 7'd1, 7'd1, 7'd3, -7'd1, 7'd1, -7'd2, -7'd2, 7'd3, -7'd1, -7'd1, 7'd0, 7'd3, 7'd1, 7'd0, -7'd1, -7'd2, 7'd0, 7'd1, 7'd4, 7'd4, -7'd1, -7'd2, 7'd2, 7'd2, 7'd2, -7'd2, 7'd2, -7'd1, 7'd4, 7'd2, -7'd3, 7'd2, 7'd0, 7'd2, 7'd1, -7'd2, -7'd1, -7'd2, 7'd0, -7'd2, 7'd0, -7'd1, 7'd3, -7'd2, 7'd2, 7'd0, 7'd1, 7'd0, 7'd0, 7'd2, 7'd2, -7'd1, -7'd3, 7'd0, -7'd4, -7'd3, 7'd0, -7'd1, 7'd0, -7'd2, 7'd1, 7'd0, 7'd0, -7'd3, -7'd1, -7'd1, 7'd2, 7'd1, -7'd2, 7'd4, -7'd2, 7'd1, 7'd1, 7'd2, -7'd1, 7'd3, 7'd4, -7'd3, -7'd1, 7'd0, -7'd2, -7'd1, 7'd0, 7'd3, 7'd3, 7'd0, -7'd1, 7'd0, 7'd3, 7'd2, -7'd1, 7'd0, 7'd1, 7'd0, 7'd0, -7'd2, 7'd3, 7'd2, -7'd1, -7'd1, 7'd1, 7'd1, 7'd0, 7'd2, 7'd3, -7'd2, 7'd2, -7'd2, 7'd1, -7'd1, -7'd1, -7'd2, -7'd1, -7'd2, -7'd3, 7'd4, -7'd1, 7'd4, -7'd1, 7'd1, -7'd2, -7'd1, 7'd0, -7'd2, 7'd0, -7'd1, -7'd2, 7'd1, -7'd1, 7'd0, 7'd3, 7'd0, 7'd1, -7'd5, 7'd1, 7'd2, 7'd3, 7'd0, 7'd1, -7'd2, 7'd0, 7'd0, -7'd2, 7'd0, -7'd2, 7'd4, -7'd1, 7'd1, 7'd0, 7'd2, 7'd1, 7'd0, -7'd4, -7'd1, -7'd1, -7'd3, -7'd2, 7'd3, -7'd1, 7'd2, 7'd3, -7'd2, 7'd1, 7'd3, 7'd2, -7'd1, 7'd1, -7'd1, -7'd1, 7'd1, -7'd1, 7'd0, 7'd2, -7'd2, 7'd0, 7'd0, 7'd1, 7'd0, -7'd1, 7'd0, 7'd0, -7'd2, 7'd1, -7'd1, 7'd0, 7'd4, -7'd2, 7'd4, 7'd2, 7'd2, 7'd1, 7'd1, -7'd2, 7'd1, 7'd1, -7'd4, -7'd2, 7'd1, 7'd0, -7'd2, 7'd3, -7'd2, -7'd2, -7'd1, 7'd1, 7'd0, -7'd2, 7'd1, -7'd4, -7'd4, 7'd0, -7'd1, -7'd4, 7'd0, 7'd2, 7'd1, 7'd3, -7'd1, 7'd1, 7'd0, 7'd4, 7'd2, -7'd3, -7'd3, -7'd1, 7'd1, -7'd3, -7'd1, -7'd1, -7'd2, 7'd0, 7'd0, 7'd2, 7'd2, 7'd4, 7'd0, -7'd3, 7'd2, -7'd4, 7'd1, 7'd3, 7'd0, 7'd0, -7'd1, 7'd1, 7'd3, -7'd2, -7'd1, 7'd2, 7'd3, 7'd0, -7'd1, -7'd2, 7'd1, -7'd1, 7'd3, -7'd2, 7'd2, -7'd1, -7'd2, 7'd3, -7'd1, 7'd0, 7'd3, -7'd2, -7'd1, 7'd0, -7'd3, -7'd1, 7'd0, -7'd2, -7'd1, -7'd1, 7'd3, 7'd0, 7'd1, -7'd2, 7'd0, 7'd2, -7'd4, 7'd2, 7'd1, 7'd4, -7'd2, 7'd1, 7'd4, 7'd1, -7'd1, 7'd1, 7'd0, -7'd1, -7'd1, -7'd4, 7'd1, -7'd3, 7'd3, 7'd2, 7'd0, 7'd2, 7'd1, 7'd3, -7'd1, -7'd1, 7'd3, 7'd4, 7'd4, 7'd0, -7'd3, -7'd2, 7'd0, 7'd2, 7'd0, -7'd2, 7'd3, 7'd1, 7'd2, -7'd3, 7'd1, -7'd2, -7'd1, 7'd2, -7'd2, 7'd0, 7'd2, 7'd1, -7'd4, -7'd3, -7'd2, -7'd4, 7'd0, -7'd3, -7'd2, 7'd2, 7'd0, 7'd2, 7'd0, -7'd1, 7'd0, 7'd1, 7'd0, 7'd1, -7'd3, 7'd0, 7'd0, -7'd4, -7'd4, -7'd3, -7'd1, -7'd2, 7'd2, -7'd1, 7'd2, -7'd4, 7'd0, -7'd1, 7'd4, 7'd1, 7'd3, 7'd1, 7'd2, 7'd1, 7'd0, -7'd4, -7'd3, 7'd0, 7'd4, -7'd1, 7'd2, -7'd1, 7'd2, 7'd2, 7'd2, 7'd2, -7'd2, -7'd1, 7'd0, 7'd0, -7'd2, 7'd1, 7'd3, -7'd1, -7'd1, 7'd1, 7'd0, 7'd0, 7'd0, -7'd3, 7'd2, 7'd2, 7'd4, 7'd1, -7'd3, -7'd2, 7'd1, 7'd0, 7'd0, -7'd4, 7'd1, -7'd1, -7'd4, 7'd3, 7'd0, -7'd4, 7'd4, 7'd3, -7'd1, 7'd2, -7'd2, 7'd2, 7'd2, -7'd3, 7'd0, -7'd3, 7'd0, 7'd3, -7'd2, -7'd1, 7'd4, 7'd1, 7'd1, 7'd1, 7'd1, -7'd1, 7'd3, 7'd3, 7'd0, 7'd1, -7'd2, -7'd1, 7'd0, -7'd4, 7'd1, -7'd2, 7'd3, -7'd4, -7'd1, -7'd2, -7'd2, 7'd4, 7'd0, 7'd0, 7'd2, -7'd2, 7'd0, -7'd1, -7'd3, -7'd2, 7'd0, 7'd1, -7'd3, 7'd1, 7'd1, -7'd1, 7'd2, 7'd0, 7'd0, 7'd1, -7'd2, -7'd2, 7'd0, 7'd3, 7'd1, -7'd2, 7'd3, 7'd2, -7'd1, 7'd2, 7'd1, -7'd3, -7'd3, -7'd2, -7'd3, 7'd0, -7'd1, 7'd2, 7'd3, 7'd3, 7'd1, -7'd1, 7'd1, -7'd4, -7'd2, 7'd1, -7'd2, 7'd3, -7'd1, -7'd3, 7'd1, 7'd1, 7'd0, -7'd1, -7'd4, 7'd0, 7'd4, -7'd2, 7'd4, 7'd1, 7'd2, 7'd1, 7'd2, -7'd2, 7'd1, 7'd2, -7'd1, -7'd1, -7'd1, -7'd4, -7'd1, 7'd3, 7'd2, -7'd3, -7'd2, -7'd2, 7'd2, -7'd1, -7'd1, -7'd3, -7'd1, 7'd2, -7'd2, -7'd3, 7'd3, -7'd1, -7'd1, -7'd1, 7'd0, -7'd2, 7'd3, -7'd3, -7'd3, 7'd0, 7'd0, -7'd2, -7'd3, -7'd2, -7'd1, 7'd3, -7'd2, 7'd2, -7'd5, -7'd2, 7'd0, -7'd2, -7'd1, 7'd0, -7'd1, 7'd1, -7'd1, 7'd0, -7'd4, 7'd0, -7'd2, 7'd2, 7'd1, 7'd1, 7'd1, -7'd3, 7'd1, -7'd1, -7'd2, 7'd1, 7'd1, 7'd0, -7'd1, 7'd1, 7'd2, -7'd1, 7'd0, 7'd0, 7'd2, 7'd3, 7'd0, -7'd1, -7'd4, 7'd2, -7'd3, 7'd2, 7'd0, -7'd3, -7'd3, 7'd2, 7'd3, 7'd1, -7'd2, 7'd0, -7'd2, 7'd0, -7'd1, -7'd1, 7'd3, -7'd2, 7'd3, 7'd2, 7'd0, 7'd3, 7'd2, 7'd0, -7'd1, 7'd0, -7'd1, 7'd3, 7'd0, 7'd4, 7'd0, 7'd2, 7'd4, -7'd1, -7'd2, 7'd0, 7'd3, 7'd3, 7'd0, -7'd1, -7'd1, 7'd0, 7'd3, -7'd3, 7'd1, 7'd0, 7'd2, 7'd1, 7'd0, 7'd1, -7'd2, 7'd2, 7'd0, 7'd3, 7'd0, 7'd2, -7'd4, 7'd2, 7'd0, -7'd2, -7'd1, 7'd0, -7'd1, 7'd1, -7'd4, 7'd2, 7'd3, -7'd1, -7'd1, 7'd1, 7'd1, -7'd2, -7'd1, 7'd1, -7'd2, -7'd2, -7'd3, -7'd2, -7'd4, 7'd0, 7'd0, 7'd2, 7'd0, -7'd1, 7'd2, -7'd1, 7'd1, 7'd2, 7'd3, 7'd3, -7'd3, -7'd1, -7'd1, 7'd4, -7'd3, 7'd2, 7'd0, 7'd0, -7'd1, -7'd1, -7'd3, -7'd3, 7'd0, 7'd0, -7'd3, -7'd3, 7'd3, 7'd0, 7'd1, 7'd2, -7'd1, 7'd1, -7'd2, 7'd1, 7'd4, 7'd4, -7'd2, 7'd2, 7'd1, 7'd2, -7'd3, 7'd4, -7'd1, -7'd3, 7'd3, -7'd3, -7'd4, -7'd2, 7'd0, -7'd2, -7'd1, 7'd4, -7'd2, -7'd2, 7'd2, 7'd2, -7'd1, 7'd2, -7'd3, 7'd0, -7'd3, -7'd3, 7'd0, -7'd2, -7'd2, 7'd0, -7'd1, -7'd1, 7'd1, 7'd1, -7'd2, 7'd1, 7'd2, 7'd1, -7'd1, -7'd2, 7'd1, -7'd1, 7'd2, 7'd4, 7'd0, 7'd2, -7'd1, 7'd0, 7'd3, -7'd2, 7'd1, 7'd1, -7'd3, -7'd1, 7'd1, 7'd1, 7'd1, 7'd1, -7'd4, -7'd3, 7'd1, 7'd1, -7'd1, 7'd1, -7'd2, 7'd1, -7'd2, 7'd4, -7'd2, 7'd1, 7'd1, 7'd1, -7'd1, -7'd3, 7'd2, -7'd1, 7'd0, 7'd3, 7'd1, 7'd3, -7'd3, -7'd3, -7'd1, 7'd0, -7'd4, 7'd3, 7'd1, 7'd0, 7'd1, -7'd2, -7'd2, -7'd2, -7'd1, 7'd1, -7'd1, -7'd2, 7'd0, 7'd2, -7'd4, 7'd4, -7'd1, -7'd4, 7'd1, -7'd1, 7'd2, 7'd2, 7'd2, -7'd1, 7'd0, 7'd0, -7'd1, 7'd4, -7'd3, -7'd3, -7'd2, 7'd3, 7'd3, -7'd1, -7'd2, 7'd1, -7'd1, 7'd2, -7'd2, -7'd2, 7'd0, 7'd1, 7'd0, 7'd1, 7'd1, -7'd1, -7'd3, -7'd2, 7'd4, 7'd3, 7'd0, 7'd3, 7'd0, -7'd4, 7'd1, 7'd2, 7'd1, 7'd0, 7'd0, 7'd4, 7'd0, -7'd1, -7'd1, -7'd1, 7'd0, 7'd3, 7'd3, -7'd1, -7'd3, -7'd2, -7'd1, -7'd3, -7'd2, 7'd1, 7'd1, -7'd1, -7'd3, 7'd1, -7'd2, -7'd3, 7'd0, 7'd4, 7'd0, -7'd3, 7'd0, -7'd3, 7'd2, 7'd0, -7'd2, -7'd1, -7'd1, 7'd1, 7'd0, 7'd1, 7'd2, -7'd4, 7'd0, 7'd3, 7'd0, -7'd1, 7'd1, 7'd0, -7'd2, -7'd2, -7'd1, -7'd2, 7'd2, -7'd2, -7'd3, 7'd0, 7'd1, 7'd1, 7'd0, -7'd4, -7'd1, -7'd2, 7'd1, -7'd1, 7'd3, 7'd4, 7'd1, -7'd4, 7'd1, 7'd4, 7'd2, -7'd2, 7'd4, 7'd0, 7'd0, 7'd2, 7'd0, -7'd3, -7'd2, 7'd0, 7'd0, -7'd4, 7'd2, 7'd2, -7'd1, 7'd3, 7'd1, 7'd1, 7'd3, 7'd4, -7'd3, 7'd0, 7'd2, -7'd2, -7'd2, 7'd0, -7'd1, 7'd0, -7'd3, -7'd1, -7'd2, -7'd1, -7'd2, 7'd2, 7'd2, -7'd4, 7'd2, 7'd3, 7'd0, -7'd2, 7'd1, 7'd1, -7'd3, -7'd2, 7'd2, -7'd2, -7'd1, 7'd1, 7'd3, -7'd2, 7'd0, 7'd4, 7'd4, 7'd2, -7'd1, -7'd1, 7'd2, 7'd0, 7'd2, 7'd2, 7'd0, -7'd2, 7'd3, 7'd2, 7'd1, -7'd4, -7'd1, -7'd4, -7'd1, 7'd3, -7'd2, 7'd1, -7'd3, -7'd2, 7'd1, 7'd0, -7'd2, -7'd1, -7'd1, 7'd0, -7'd2, 7'd1, 7'd0, -7'd2, 7'd1, 7'd0, 7'd3, 7'd1, 7'd1, 7'd0, 7'd1, -7'd2, -7'd4, 7'd1, 7'd0, -7'd1, -7'd4, 7'd0, 7'd2, 7'd2, 7'd1, 7'd1, 7'd1, -7'd1, -7'd1, 7'd4, 7'd0, -7'd2, -7'd2, 7'd1, -7'd3, 7'd1, 7'd2, 7'd0, -7'd2, -7'd1, 7'd1, -7'd1, -7'd5, -7'd2, -7'd2, -7'd3, -7'd3, 7'd1, 7'd1, -7'd1, 7'd3, -7'd1, 7'd3, -7'd1, 7'd4, 7'd1, -7'd1, 7'd1, 7'd1, -7'd2, 7'd1, -7'd3, 7'd0, 7'd2, 7'd2, 7'd0, -7'd3, -7'd4, 7'd0, 7'd3, -7'd2, -7'd1, -7'd1, 7'd2, 7'd2, -7'd3, -7'd2, -7'd1, -7'd1, -7'd2, -7'd1, 7'd1, 7'd1, -7'd1, -7'd4, 7'd1, -7'd1, 7'd1, 7'd3, 7'd0, 7'd0, 7'd1, -7'd1, 7'd0, 7'd0, -7'd3, -7'd2, 7'd0, -7'd2, 7'd1, -7'd1, -7'd3, 7'd2, -7'd1, -7'd1, -7'd1, 7'd0, 7'd3, -7'd2, 7'd2, -7'd2, 7'd0, 7'd2, 7'd2, -7'd1, -7'd1, 7'd0, -7'd3, -7'd2, 7'd1, -7'd1, -7'd2, 7'd1, -7'd1, 7'd2, 7'd4, 7'd0, 7'd0, 7'd1, 7'd3, 7'd1, 7'd1, 7'd0, 7'd0, -7'd2, 7'd2, 7'd3, -7'd4, 7'd3, 7'd0, -7'd1, 7'd2, 7'd2, 7'd2, 7'd2, 7'd2, -7'd4, -7'd1, -7'd2, -7'd3, -7'd2, -7'd1, 7'd3, 7'd0, 7'd3, -7'd1, 7'd1, 7'd4, 7'd1, -7'd4, -7'd2, 7'd0, 7'd2, 7'd0, -7'd4, -7'd2, -7'd1, 7'd3, 7'd2, 7'd0, 7'd1, 7'd1, -7'd1, -7'd3, 7'd1, -7'd2, 7'd3, 7'd1, -7'd3, 7'd1, -7'd1, -7'd1, -7'd1, 7'd0, 7'd0, -7'd3, -7'd2, 7'd0, -7'd4, -7'd2, 7'd3, -7'd2, 7'd0, 7'd2, -7'd1, 7'd3, -7'd1, -7'd4, -7'd2, -7'd1, 7'd0, -7'd2, -7'd2, 7'd4, 7'd4, 7'd2, -7'd1, 7'd0, -7'd1, 7'd2, 7'd2, -7'd3, -7'd3, 7'd1, 7'd1, 7'd0, -7'd1, 7'd2, -7'd2, -7'd1, 7'd1, -7'd1, -7'd3, -7'd1, -7'd5, 7'd2, 7'd2, -7'd3, -7'd3, -7'd1, -7'd1, -7'd2, 7'd2, 7'd0, 7'd3, 7'd2, 7'd2, -7'd1, -7'd1, 7'd1, 7'd2, 7'd2, -7'd1, -7'd1, 7'd1, -7'd1, -7'd2, -7'd4, -7'd1, 7'd1, 7'd4, 7'd2, 7'd1, 7'd1, -7'd1, 7'd1, 7'd2, -7'd4, -7'd1, 7'd2, 7'd2, -7'd1, 7'd0, 7'd0, 7'd0, 7'd1, 7'd3, 7'd2, 7'd1, -7'd1, -7'd1, 7'd2, 7'd2, 7'd2, 7'd3, -7'd2, 7'd3, -7'd1, 7'd1, 7'd3, 7'd2, 7'd1, -7'd3, 7'd0, -7'd1, -7'd1, 7'd0, 7'd1, 7'd0, 7'd0, 7'd3, -7'd3, -7'd1, -7'd2, -7'd1, -7'd4, 7'd1, 7'd3, 7'd1, 7'd0, 7'd0, 7'd1, -7'd3, 7'd1, -7'd4, 7'd0, 7'd1, 7'd1, 7'd1, -7'd2, 7'd0, 7'd3, 7'd0, 7'd4, -7'd2, -7'd1, -7'd1, -7'd1, -7'd1, 7'd2, -7'd1, -7'd1, 7'd0, 7'd1, 7'd0, 7'd1, 7'd2, -7'd1, -7'd1, 7'd1, 7'd4, 7'd2, -7'd4, 7'd1, 7'd0, 7'd2, -7'd1, 7'd2, -7'd3, 7'd3, 7'd0, 7'd3, -7'd1, -7'd3, 7'd1, -7'd1, -7'd2, -7'd3, -7'd2, 7'd0, 7'd0, -7'd2, 7'd2, 7'd0, 7'd4, 7'd2, 7'd0, -7'd3, -7'd2, -7'd2, 7'd0, -7'd2, 7'd3, -7'd2, -7'd1, 7'd4, -7'd1, 7'd0, -7'd4, -7'd2, 7'd3, -7'd3, 7'd0, -7'd1, -7'd3, -7'd3, 7'd0, 7'd2, 7'd1, 7'd1, -7'd3, 7'd0, 7'd3, -7'd2, 7'd1, 7'd2, 7'd0, 7'd3, -7'd3, 7'd0, 7'd0, -7'd3, 7'd2, 7'd1, -7'd4, 7'd0, 7'd1, -7'd2, -7'd3, 7'd1, 7'd1, -7'd2, 7'd1, 7'd2, 7'd1, 7'd1, 7'd4, -7'd1, 7'd2, -7'd3, -7'd3, 7'd3, -7'd1, 7'd1, 7'd0, 7'd3, -7'd3, 7'd1, 7'd2, 7'd3, 7'd1, -7'd1, 7'd3, 7'd3, 7'd3, -7'd4, 7'd0, 7'd0, 7'd2, 7'd4, 7'd5, 7'd2, -7'd2, -7'd2, 7'd0, 7'd0, 7'd0, 7'd0, -7'd1, 7'd1, 7'd4, 7'd1, -7'd1, 7'd0, -7'd1, -7'd3, 7'd0, 7'd2, 7'd2, -7'd2, -7'd1, -7'd2, 7'd0, 7'd1, 7'd3, -7'd2, 7'd3, 7'd0, 7'd0, 7'd0, -7'd2, 7'd3, 7'd1, -7'd3, 7'd0, -7'd3, 7'd0, 7'd2, -7'd3, -7'd2, 7'd3, 7'd4, 7'd2, 7'd1, 7'd0, -7'd3, -7'd1, -7'd2, 7'd3, -7'd3, -7'd1, -7'd3, 7'd2, 7'd2, -7'd4, 7'd1, 7'd0, -7'd1, -7'd1, -7'd2, -7'd3, 7'd1, 7'd2, -7'd1, 7'd2, 7'd0, 7'd1, -7'd1, 7'd3, 7'd1, 7'd2, -7'd2, 7'd2, -7'd3, -7'd1, -7'd4, 7'd0, 7'd1, -7'd3, 7'd4, 7'd1, -7'd3, -7'd1, -7'd1, 7'd3, -7'd1, 7'd0, 7'd1, 7'd3, -7'd1, 7'd1, 7'd2, 7'd2, 7'd3, 7'd0, 7'd1, 7'd4, 7'd1, -7'd1, 7'd1, 7'd1, -7'd1, 7'd4, -7'd4, -7'd2, 7'd4, -7'd1, 7'd1, 7'd1, -7'd1, -7'd1, 7'd2, 7'd3, 7'd2, -7'd1, 7'd3, -7'd2, 7'd0, -7'd1, 7'd0, 7'd0, 7'd1, -7'd3, 7'd0, -7'd2, -7'd2, -7'd3, -7'd4, 7'd1, -7'd2, 7'd0, -7'd1, -7'd1, 7'd1, -7'd1, 7'd3, 7'd1, -7'd2, 7'd2, -7'd1, -7'd1, 7'd0, 7'd2, -7'd2, -7'd3, 7'd0, 7'd0, 7'd0, -7'd2, -7'd4, 7'd1, 7'd2, 7'd1, -7'd2, -7'd1, 7'd0, 7'd0, 7'd4, 7'd0, 7'd0, 7'd3, 7'd2, 7'd3, -7'd1, 7'd0, -7'd1, -7'd2, -7'd2, 7'd2, -7'd2, -7'd2, 7'd3, -7'd1, -7'd2, -7'd1, 7'd1, -7'd3, 7'd2, 7'd3, -7'd1, 7'd1, -7'd3, 7'd2, 7'd0, -7'd1, 7'd0, -7'd2, 7'd2, 7'd0, 7'd1, -7'd1, -7'd1, 7'd1, -7'd4, -7'd2, 7'd0, 7'd1, -7'd2, 7'd3, 7'd4, 7'd3, 7'd0, -7'd2, 7'd3, 7'd3, 7'd2, -7'd4, -7'd3, 7'd2, 7'd0, 7'd3, 7'd2, 7'd0, 7'd2, 7'd0, 7'd0, -7'd1, -7'd4, 7'd4, 7'd3, 7'd1, -7'd3, 7'd0, -7'd1, -7'd3, 7'd2, -7'd2, -7'd4, -7'd1, 7'd1, -7'd3, 7'd0, 7'd1, 7'd4, 7'd1, 7'd2, 7'd0, 7'd3, 7'd3, 7'd4, -7'd1, 7'd1, -7'd1, 7'd2, 7'd5, -7'd1, 7'd0, 7'd1, -7'd4, 7'd3, -7'd2, 7'd0, 7'd1, 7'd4, 7'd1, 7'd2, 7'd0, 7'd1, 7'd1, 7'd0, 7'd1, -7'd1, 7'd1, 7'd0, -7'd2, 7'd1, 7'd2, 7'd0, 7'd2, 7'd2, -7'd3, -7'd4, 7'd1, 7'd0, 7'd0, 7'd0, -7'd2, 7'd3, -7'd1, -7'd1, -7'd3, -7'd1, -7'd3, -7'd3, 7'd4, -7'd2, -7'd2, -7'd2, -7'd1, 7'd2, 7'd0, 7'd4, -7'd1, -7'd1, 7'd0, 7'd0, 7'd3, -7'd4, 7'd0, 7'd2, 7'd4, -7'd1, -7'd1, 7'd0, -7'd1, -7'd4, -7'd1, -7'd3, -7'd2, 7'd1, -7'd2, 7'd1, -7'd3, 7'd0, -7'd2, 7'd1, 7'd2, 7'd2, 7'd5, -7'd2, 7'd2, 7'd1, -7'd4, 7'd2, 7'd1, -7'd1, 7'd0, 7'd1, 7'd1, 7'd0, 7'd1, -7'd2, -7'd4, 7'd2, 7'd0, 7'd3, -7'd1, -7'd3, -7'd2, -7'd2, 7'd2, 7'd1, -7'd2, -7'd1, 7'd0, 7'd2, 7'd0, -7'd2, -7'd1, 7'd3, -7'd2, 7'd0, -7'd1, 7'd2, 7'd1, 7'd2, -7'd1, 7'd1, -7'd1, -7'd1, -7'd2, -7'd3, 7'd1, -7'd1, 7'd0, 7'd0, 7'd1, 7'd3, 7'd0, 7'd2, 7'd0, -7'd1, 7'd4, 7'd1, 7'd0, 7'd0, 7'd0, -7'd3, -7'd3, 7'd2, -7'd2, 7'd0, 7'd1, 7'd1, -7'd2, 7'd4, -7'd1, -7'd2, 7'd3, 7'd0, -7'd2, 7'd0, 7'd2, 7'd2, -7'd3, -7'd2, 7'd1, 7'd2, 7'd0, 7'd2, 7'd0, 7'd0, -7'd2, -7'd1, 7'd2, -7'd2, 7'd3, 7'd0, 7'd3, 7'd1, 7'd2, -7'd1, -7'd3, -7'd1, 7'd0, -7'd2, 7'd0, 7'd1, 7'd2, -7'd2, 7'd4, -7'd1, -7'd1, -7'd1, 7'd4, 7'd2, 7'd0, 7'd0, 7'd1, 7'd1, 7'd1, 7'd0, 7'd4, -7'd3, 7'd3, 7'd0, 7'd3, 7'd1, 7'd4, -7'd2, 7'd1, 7'd1, -7'd3, -7'd1, 7'd2, 7'd1, -7'd2, -7'd2, -7'd2, 7'd0, 7'd1, 7'd0, 7'd1, 7'd1, -7'd2, 7'd0, -7'd4, 7'd1, -7'd3, 7'd1, -7'd1, -7'd1, 7'd1, -7'd2, -7'd1, -7'd3, 7'd1, 7'd3, -7'd1, 7'd0, -7'd3, -7'd4, 7'd0, 7'd1, -7'd1, 7'd1, -7'd1, 7'd2, 7'd3, 7'd4, 7'd2, 7'd3, -7'd3, -7'd2, -7'd1, 7'd0, -7'd3, 7'd4, -7'd2, -7'd1, -7'd2, 7'd0, -7'd1, -7'd1, 7'd0, -7'd3, -7'd1, 7'd0, 7'd0, -7'd3, 7'd0, -7'd3, -7'd1, -7'd1, -7'd2, 7'd1, 7'd1, -7'd1, -7'd3, 7'd2, 7'd0, 7'd0, -7'd2, 7'd0, -7'd2, 7'd0, -7'd2, 7'd2, -7'd3, -7'd1, -7'd4, 7'd1, 7'd1, 7'd0, 7'd1, 7'd1, -7'd1, 7'd3, 7'd4, -7'd4, 7'd0, -7'd4, 7'd2, 7'd0, 7'd4, 7'd1, -7'd1, 7'd1, 7'd1, -7'd1, -7'd2, 7'd1, -7'd2, 7'd4, 7'd1, -7'd2, 7'd0, -7'd1, -7'd2, -7'd1, 7'd2, 7'd0, -7'd1, -7'd2, -7'd1, -7'd1, -7'd2, 7'd1, 7'd2, 7'd0, 7'd1, 7'd0, -7'd1, 7'd1, -7'd2, -7'd1, -7'd3, 7'd0, -7'd4, -7'd2, -7'd1, -7'd2, 7'd0, 7'd3, 7'd2, 7'd1, 7'd3, -7'd1, 7'd1, -7'd3, -7'd1, -7'd1, -7'd1, -7'd1, 7'd2, 7'd0, 7'd3, 7'd1, 7'd0, 7'd0, -7'd1, 7'd4, 7'd1, -7'd1, 7'd1, -7'd2, 7'd0, 7'd2, 7'd3, 7'd2, -7'd1, -7'd1, -7'd1, -7'd1, 7'd1, 7'd2, 7'd1, 7'd1, -7'd2, 7'd3, -7'd1, 7'd0, 7'd0, 7'd0, -7'd2, -7'd3, 7'd2, 7'd0, -7'd1, -7'd1, -7'd2, -7'd2, 7'd3, 7'd1, -7'd1, 7'd0, -7'd2, 7'd2, -7'd4, 7'd1, 7'd0, 7'd2, -7'd3, 7'd2, 7'd1, -7'd2, 7'd0, -7'd4, 7'd1, 7'd2, 7'd3, 7'd1, -7'd2, 7'd2, 7'd0, -7'd1, 7'd2, 7'd0, -7'd2, 7'd2, 7'd2, 7'd0, -7'd1, 7'd2, -7'd1, -7'd1, 7'd0, -7'd1, 7'd0, 7'd2, 7'd1, -7'd4, 7'd4, -7'd1, -7'd3, -7'd2, 7'd1, -7'd1, -7'd1, 7'd0, 7'd2, -7'd2, 7'd1, 7'd1, 7'd2, 7'd2, -7'd1, -7'd2, -7'd1, 7'd1, 7'd2, 7'd1, 7'd0, -7'd3, 7'd3, 7'd0, 7'd3, -7'd1, 7'd0, -7'd2, 7'd2, -7'd3, 7'd0, 7'd0, -7'd2, 7'd3, 7'd0, -7'd3, 7'd1, 7'd0, 7'd3, -7'd1, 7'd1, -7'd1, -7'd2, -7'd1, 7'd0, 7'd1, 7'd3, -7'd5, -7'd1, -7'd1, 7'd2, 7'd4, -7'd2, -7'd1, 7'd3, 7'd2, 7'd2, -7'd2, 7'd3, -7'd1, -7'd1, 7'd1, 7'd0, -7'd1, 7'd0, -7'd2, 7'd3, -7'd2, 7'd4, -7'd2, -7'd2, -7'd1, 7'd3, 7'd3, 7'd2, 7'd0, 7'd0, 7'd2, -7'd2, -7'd1, -7'd4, 7'd1, 7'd0, 7'd0, 7'd4, 7'd4, 7'd1, 7'd1, 7'd3, 7'd1, 7'd3, -7'd1, 7'd1, 7'd0, -7'd3, 7'd3, -7'd2, 7'd4, -7'd1, -7'd4, 7'd1, 7'd3, 7'd0, 7'd0, 7'd0, 7'd1, -7'd1, -7'd3, -7'd4, 7'd3, -7'd4, -7'd3, -7'd3, 7'd1, -7'd1, -7'd1, 7'd0, -7'd1, -7'd3, 7'd1, 7'd0, 7'd0, 7'd2, -7'd2, 7'd1, 7'd1, -7'd3, 7'd1, 7'd2, -7'd2, 7'd0, 7'd1, 7'd1, 7'd2, -7'd1, 7'd2, 7'd1, -7'd1, -7'd3, 7'd1, 7'd3,  5'd0, 5'd0, 5'd0, 5'd0, 5'd0, 5'd0, 5'd0, 5'd0, 5'd0, 5'd0, 5'd0, 5'd0, 5'd0, 5'd0, 5'd0, 5'd0, 5'd0, 5'd0, 5'd0, 5'd0, 5'd0, 5'd0, 5'd0, 5'd0, 5'd0, 5'd0, 5'd0, 5'd0, 5'd0, 5'd0, 5'd0, 5'd0, 5'd2, -5'd2, 5'd2, 5'd2, -5'd2, -5'd1, 5'd0, 5'd1, -5'd2, 5'd0, -5'd1, 5'd2, 5'd1, 5'd0, 5'd0, 5'd4, 5'd3, 5'd1, 5'd0, 5'd1, 5'd0, -5'd2, -5'd4, -5'd4, 5'd3, 5'd0, 5'd0, -5'd2, -5'd1, 5'd1, -5'd2, 5'd3, 5'd5, -5'd3, -5'd1, 5'd3, 5'd1, 5'd0, 5'd0, -5'd1, 5'd4, -5'd1, -5'd1, -5'd2, -5'd4, 5'd1, -5'd5, 5'd1, 5'd4, -5'd1, 5'd2, -5'd1, -5'd1, 5'd0, 5'd1, -5'd1, 5'd0, -5'd4, -5'd2, 5'd4, 5'd4, -5'd4, -5'd3, -5'd2, 5'd1, 5'd1, -5'd4, -5'd3, -5'd1, -5'd2, -5'd4, -5'd1, 5'd4, -5'd4, 5'd0, -5'd1, -5'd1, -5'd1, 5'd1, 5'd0, 5'd0, 5'd0, -5'd5, -5'd4, 5'd1, -5'd4, -5'd1, 5'd1, 5'd1, 5'd0, -5'd1, 5'd2, -5'd4, 5'd3, -5'd2, -5'd1, 5'd2, 5'd0, -5'd2, 5'd0, -5'd5, 5'd2, 5'd0, 5'd0, 5'd2, 5'd3, 5'd3, 5'd1, -5'd1, 5'd3, -5'd4, -5'd2, 5'd3, 5'd5, 5'd4, -5'd3, -5'd2, -5'd2, -5'd1, 5'd1, 5'd0, 5'd1, 5'd0, -5'd1, 5'd3, -5'd3, 5'd3, -5'd2, -5'd3, 5'd2, -5'd2, -5'd3, 5'd1, 5'd2, -5'd2, 5'd0, 5'd0, -5'd2, 5'd1, 5'd1, 5'd0, 5'd0, 5'd4, 5'd2, -5'd1, -5'd1, 5'd2, 5'd1, -5'd4, 5'd2, 5'd0, -5'd2, 5'd3, 5'd2, 5'd1, 5'd0, 5'd0, 5'd2, 5'd1, -5'd3, -5'd1, -5'd2, 5'd2, -5'd3, -5'd3, -5'd1, -5'd4, 5'd0, -5'd2, -5'd2, 5'd1, 5'd0, 5'd1, 5'd5, -5'd5, 5'd3, -5'd1, -5'd5, 5'd4, 5'd1, 5'd3, 5'd0, 5'd1, -5'd1, -5'd2, -5'd4, 5'd4, -5'd2, 5'd1, -5'd1, -5'd1, 5'd0, -5'd4, 5'd4, 5'd4, -5'd1, -5'd1, 5'd1, 5'd3, -5'd2, 5'd4, 5'd1, 5'd0, 5'd0, -5'd2, -5'd2, 5'd1, -5'd1, -5'd3, 5'd1, -5'd5, -5'd1, -5'd1, 5'd2, 5'd2, 5'd1, -5'd4, -5'd2, -5'd2, -5'd2, 5'd1, -5'd1, -5'd1, -5'd2, -5'd1, -5'd1, 5'd2, -5'd1, -5'd4, 5'd3, 5'd0, 5'd4, 5'd1, -5'd1, 5'd0, 5'd2, -5'd2, 5'd3, 5'd2, 5'd2, 5'd0, 5'd0, 5'd3, -5'd1, -5'd1, -5'd2, 5'd0, -5'd3, 5'd3, -5'd2, 5'd2, -5'd1, 5'd3, 5'd4, -5'd2, 5'd3, 5'd1, 5'd1, -5'd1, -5'd1, -5'd1, -5'd3, -5'd1, -5'd2, 5'd0, -5'd2, -5'd4, -5'd1, 5'd1, -5'd3, -5'd2, 5'd1, 5'd2, 5'd1, -5'd1, -5'd3, -5'd1, 5'd1, 5'd0, -5'd1, -5'd4, -5'd1, 5'd1, -5'd2, -5'd1, 5'd0, 5'd0, 5'd0, -5'd3, 5'd0, -5'd1, -5'd1, -5'd2, 5'd1, 5'd2, -5'd5, 5'd4, 5'd1, 5'd2, 5'd0, 5'd0, 5'd1, 5'd0, 5'd0, 5'd1, 5'd2, 5'd0, 5'd1, 5'd3, -5'd2, -5'd2, -5'd3, -5'd2, 5'd1, 5'd2, 5'd0, 5'd3, -5'd1, 5'd3, -5'd1, 5'd3, -5'd2, 5'd1, -5'd4, 5'd1, 5'd1, -5'd1, 5'd1, -5'd5, 5'd4, 5'd2, -5'd1, 5'd0, -5'd2, -5'd2, 5'd2, 5'd1, 5'd3, 5'd3, 5'd1, -5'd3, 5'd3, -5'd1, 5'd4, -5'd3, 5'd3, -5'd5, -5'd1, -5'd1, 5'd3, 5'd0, 5'd0, 5'd0, 5'd2, 5'd0, 5'd2, 5'd2, -5'd2, -5'd1, -5'd1, -5'd2, 5'd0, 5'd0, 5'd0, 5'd3, 5'd2, 5'd2, 5'd0, 5'd1, 5'd1, 5'd0, -5'd1, -5'd3, 5'd2, -5'd1, 5'd2, 5'd4, 5'd2, 5'd2, 5'd2, 5'd0, 5'd4, -5'd2, 5'd1, -5'd3, -5'd4, -5'd2, 5'd5, 5'd1, -5'd3, -5'd2, -5'd1, -5'd5, 5'd3, 5'd0, 5'd0, 5'd2, 5'd0, 5'd0, -5'd1, 5'd1, -5'd1, 5'd3, 5'd3, 5'd4, -5'd1, 5'd1, -5'd1, -5'd1, -5'd1, -5'd1, -5'd3, 5'd1, 5'd4, 5'd3, -5'd3, 5'd2, -5'd1, 5'd0, 5'd4, 5'd0, -5'd3, -5'd1, -5'd2, 5'd3, 5'd2, -5'd1, 5'd1, -5'd1, 5'd2, -5'd1, 5'd2, 5'd0, 5'd1, 5'd1, -5'd3, -5'd1, 5'd5, 5'd4, -5'd4, 5'd1, 5'd0, 5'd2, -5'd1, 5'd1, 5'd0, -5'd4, 5'd5, 5'd3, -5'd1, -5'd2, 5'd5, 5'd0, 5'd1, -5'd3, 5'd2, 5'd2, -5'd2, 5'd1, -5'd1, -5'd2, -5'd1, 5'd3, 5'd0, -5'd1, -5'd4, -5'd3, -5'd2, 5'd2, -5'd1, -5'd2, -5'd5, -5'd2, 5'd1, 5'd1, 5'd5, 5'd0, 5'd4, 5'd5, 5'd5, 5'd1, 5'd2, 5'd2, 5'd2, 5'd2, -5'd1, 5'd0, 5'd0, 5'd3, 5'd2, -5'd2, 5'd2, 5'd0, -5'd3, -5'd2, 5'd4, 5'd1, -5'd3, -5'd1, 5'd1, 5'd0, 5'd3, 5'd1, 5'd1, 5'd1, -5'd2, -5'd1, 5'd0, -5'd2, 5'd0, -5'd2, -5'd4, 5'd0, 5'd4, 5'd2, 5'd1, -5'd2, -5'd2, 5'd0, -5'd2, -5'd3, -5'd1, 5'd1, 5'd0, -5'd1, -5'd1, -5'd1, -5'd1, -5'd1, -5'd2, 5'd4, 5'd0, 5'd2, -5'd1, 5'd1, -5'd4, 5'd1, 5'd3, 5'd3, -5'd1, 5'd2, 5'd1, 5'd0, 5'd0, 5'd1, -5'd1, 5'd2, -5'd3, 5'd3, 5'd0, -5'd3, -5'd1, 5'd3, 5'd1, -5'd2, -5'd3, 5'd2, -5'd2, 5'd1, 5'd3, -5'd4, 5'd1, 5'd1, -5'd1, 5'd2, -5'd2, 5'd2, -5'd4, 5'd1, -5'd3, 5'd2, 5'd0, 5'd0, 5'd3, -5'd4, -5'd2, 5'd2, 5'd1, -5'd2, -5'd1, 5'd2, 5'd0, -5'd2, -5'd4, 5'd0, 5'd1, -5'd1, 5'd1, 5'd0, 5'd0, 5'd1, 5'd1, 5'd0, 5'd2, 5'd3, -5'd1, -5'd1, 5'd0, -5'd1, -5'd3, 5'd0, -5'd2, 5'd2, -5'd1, 5'd2, 5'd4, -5'd1, -5'd1, -5'd1, 5'd0, 5'd4, 5'd0, -5'd3, 5'd0, 5'd4, 5'd1, -5'd2, -5'd1, 5'd1, 5'd0, -5'd5, 5'd0, -5'd1, -5'd1, -5'd2, 5'd0, -5'd3, -5'd1, 5'd2, 5'd1, 5'd4, 5'd2, 5'd1, 5'd3, 5'd2, 5'd1, 5'd1, -5'd1, 5'd0, -5'd1, 5'd0, 5'd0, -5'd3, -5'd1, -5'd3, 5'd2, 5'd5, 5'd3, -5'd3, 5'd0, 5'd3, 5'd0, 5'd0, 5'd3, 5'd3, 5'd1, 5'd1, -5'd2, 5'd3, -5'd1, 5'd4, 5'd0, -5'd2, -5'd1, 5'd2, 5'd3, -5'd1, 5'd2, -5'd2, -5'd4, -5'd3, -5'd2, 5'd3, 5'd0, 5'd3, 5'd0, -5'd3, 5'd2, -5'd3, 5'd2, 5'd5, -5'd3, 5'd4, 5'd0, -5'd3, -5'd3, -5'd1, -5'd1, -5'd2, -5'd3, 5'd1, 5'd3, 5'd1, 5'd0, 5'd2, -5'd2, 5'd2, 5'd3, -5'd3, 5'd3, -5'd2, -5'd2, 5'd1, 5'd1, -5'd3, -5'd1, 5'd0, -5'd1, -5'd4, 5'd3, -5'd5, 5'd1, 5'd1, -5'd1, 5'd0, -5'd2, 5'd0, 5'd2, 5'd3, 5'd0, 5'd2, 5'd0, -5'd3, 5'd1, -5'd1, -5'd1, 5'd1, -5'd1, 5'd2, 5'd0, 5'd4, -5'd1, -5'd2, 5'd2, 5'd4, 5'd1, -5'd2, -5'd4, -5'd2, 5'd3, -5'd5, -5'd3, -5'd2, 5'd2, -5'd1, 5'd4, -5'd2, 5'd3, -5'd1, -5'd1, -5'd2, 5'd3, -5'd2, 5'd2, -5'd1, 5'd4, 5'd2, 5'd2, 5'd0, 5'd4, 5'd1, -5'd1, 5'd0, 5'd2, 5'd1, -5'd2, 5'd1, 5'd1, -5'd4, 5'd0, -5'd1, 5'd1, -5'd3, 5'd4, 5'd4, 5'd0, 5'd3, 5'd0, -5'd3, 5'd0, 5'd0, -5'd1, 5'd2, -5'd2, 5'd1, 5'd0, -5'd3, 5'd1, -5'd2, -5'd2, 5'd1, -5'd1, -5'd2, 5'd1, -5'd1, 5'd1, 5'd1, 5'd1, -5'd1, 5'd3 };

  logic clk=0, rstn=1, copy=0, k=0;
  logic [XD-1:0][XB-1:0] x;
  logic [YD-1:0][YB-1:0] y;

  model model (.*);

  initial forever #5ns clk = !clk;

  int fd, status;
  localparam DIR = "D:/research/tritonRTL/test/vectors/";
  initial begin
    fd = $fopen({DIR,"x.txt"}, "r");
    for (int xn=0; xn<XD; xn++)
      status = $fscanf(fd, "%d", x[xn]);
    $fclose(fd);

    @(posedge clk) #1ns;
    
    for (int i=0; i<WEIGHTS_B; i++) begin
      k <= weights[i];
      copy <= 1;
      @(posedge clk) #1ns;
    end
    copy = 0;

    @(posedge clk);

    fd = $fopen({DIR,"y6_sim.txt"}, "w");
    for (int yn=0; yn<YD; yn++)
      $fdisplay(fd, "%d", model.act6_y[yn]);
    $fclose(fd);

    $finish();
  end
endmodule